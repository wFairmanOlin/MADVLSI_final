magic
tech sky130A
timestamp 1620673627
<< xpolycontact >>
rect 0 1970 35 2190
rect 0 0 35 220
rect 160 1970 195 2190
rect 160 0 195 220
rect 320 1970 355 2190
rect 320 0 355 220
rect 480 1970 515 2190
rect 480 0 515 220
rect 640 1970 675 2190
rect 640 0 675 220
rect 800 1970 835 2190
rect 800 0 835 220
rect 960 1970 995 2190
rect 960 0 995 220
rect 1120 1970 1155 2190
rect 1120 0 1155 220
rect 1280 1970 1315 2190
rect 1280 0 1315 220
rect 1440 1970 1475 2190
rect 1440 0 1475 220
<< xpolyres >>
rect 0 220 35 1970
rect 160 220 195 1970
rect 320 220 355 1970
rect 480 220 515 1970
rect 640 220 675 1970
rect 800 220 835 1970
rect 960 220 995 1970
rect 1120 220 1155 1970
rect 1280 220 1315 1970
rect 1440 220 1475 1970
<< locali >>
rect 35 1970 160 2190
rect 355 1970 480 2190
rect 675 1970 800 2190
rect 995 1970 1120 2190
rect 1315 1970 1440 2190
rect 195 0 320 220
rect 515 0 640 220
rect 835 0 960 220
rect 1155 0 1280 220
<< end >>
