magic
tech sky130A
timestamp 1620622228
<< nmos >>
rect 0 400 60 550
rect 110 400 170 550
rect 220 400 280 550
rect 330 400 390 550
rect 440 400 500 550
rect 550 400 610 550
rect 660 400 720 550
rect 770 400 830 550
rect 880 400 940 550
rect 990 400 1050 550
rect 1100 400 1160 550
rect 1210 400 1270 550
rect 1320 400 1380 550
rect 0 0 60 150
rect 110 0 170 150
rect 220 0 280 150
rect 330 0 390 150
rect 440 0 500 150
rect 550 0 610 150
rect 660 0 720 150
rect 770 0 830 150
rect 880 0 940 150
rect 990 0 1050 150
rect 1100 0 1160 150
rect 1210 0 1270 150
rect 1320 0 1380 150
<< ndiff >>
rect -50 535 0 550
rect -50 415 -35 535
rect -15 415 0 535
rect -50 400 0 415
rect 60 535 110 550
rect 60 415 75 535
rect 95 415 110 535
rect 60 400 110 415
rect 170 535 220 550
rect 170 415 185 535
rect 205 415 220 535
rect 170 400 220 415
rect 280 535 330 550
rect 280 415 295 535
rect 315 415 330 535
rect 280 400 330 415
rect 390 535 440 550
rect 390 415 405 535
rect 425 415 440 535
rect 390 400 440 415
rect 500 535 550 550
rect 500 415 515 535
rect 535 415 550 535
rect 500 400 550 415
rect 610 535 660 550
rect 610 415 625 535
rect 645 415 660 535
rect 610 400 660 415
rect 720 535 770 550
rect 720 415 735 535
rect 755 415 770 535
rect 720 400 770 415
rect 830 400 880 550
rect 940 535 990 550
rect 940 415 955 535
rect 975 415 990 535
rect 940 400 990 415
rect 1050 535 1100 550
rect 1050 415 1065 535
rect 1085 415 1100 535
rect 1050 400 1100 415
rect 1160 535 1210 550
rect 1160 415 1175 535
rect 1195 415 1210 535
rect 1160 400 1210 415
rect 1270 535 1320 550
rect 1270 415 1285 535
rect 1305 415 1320 535
rect 1270 400 1320 415
rect 1380 535 1430 550
rect 1380 415 1395 535
rect 1415 415 1430 535
rect 1380 400 1430 415
rect -50 135 0 150
rect -50 15 -35 135
rect -15 15 0 135
rect -50 0 0 15
rect 60 135 110 150
rect 60 15 75 135
rect 95 15 110 135
rect 60 0 110 15
rect 170 135 220 150
rect 170 15 185 135
rect 205 15 220 135
rect 170 0 220 15
rect 280 135 330 150
rect 280 15 295 135
rect 315 15 330 135
rect 280 0 330 15
rect 390 135 440 150
rect 390 15 405 135
rect 425 15 440 135
rect 390 0 440 15
rect 500 135 550 150
rect 500 15 515 135
rect 535 15 550 135
rect 500 0 550 15
rect 610 135 660 150
rect 610 15 625 135
rect 645 15 660 135
rect 610 0 660 15
rect 720 135 770 150
rect 720 15 735 135
rect 755 15 770 135
rect 720 0 770 15
rect 830 0 880 150
rect 940 135 990 150
rect 940 15 955 135
rect 975 15 990 135
rect 940 0 990 15
rect 1050 135 1100 150
rect 1050 15 1065 135
rect 1085 15 1100 135
rect 1050 0 1100 15
rect 1160 135 1210 150
rect 1160 15 1175 135
rect 1195 15 1210 135
rect 1160 0 1210 15
rect 1270 135 1320 150
rect 1270 15 1285 135
rect 1305 15 1320 135
rect 1270 0 1320 15
rect 1380 135 1430 150
rect 1380 15 1395 135
rect 1415 15 1430 135
rect 1380 0 1430 15
<< ndiffc >>
rect -35 415 -15 535
rect 75 415 95 535
rect 185 415 205 535
rect 295 415 315 535
rect 405 415 425 535
rect 515 415 535 535
rect 625 415 645 535
rect 735 415 755 535
rect 955 415 975 535
rect 1065 415 1085 535
rect 1175 415 1195 535
rect 1285 415 1305 535
rect 1395 415 1415 535
rect -35 15 -15 135
rect 75 15 95 135
rect 185 15 205 135
rect 295 15 315 135
rect 405 15 425 135
rect 515 15 535 135
rect 625 15 645 135
rect 735 15 755 135
rect 955 15 975 135
rect 1065 15 1085 135
rect 1175 15 1195 135
rect 1285 15 1305 135
rect 1395 15 1415 135
<< psubdiff >>
rect -100 535 -50 550
rect -100 415 -85 535
rect -65 415 -50 535
rect -100 400 -50 415
rect 1430 535 1480 550
rect 1430 415 1445 535
rect 1465 415 1480 535
rect 1430 400 1480 415
rect -100 135 -50 150
rect -100 15 -85 135
rect -65 15 -50 135
rect -100 0 -50 15
rect 1430 135 1480 150
rect 1430 15 1445 135
rect 1465 15 1480 135
rect 1430 0 1480 15
<< psubdiffcont >>
rect -85 415 -65 535
rect 1445 415 1465 535
rect -85 15 -65 135
rect 1445 15 1465 135
<< poly >>
rect 220 590 280 605
rect 220 570 240 590
rect 260 570 280 590
rect 0 550 60 565
rect 110 550 170 565
rect 220 550 280 570
rect 660 590 720 605
rect 660 570 680 590
rect 700 570 720 590
rect 330 550 390 565
rect 440 550 500 565
rect 550 550 610 565
rect 660 550 720 570
rect 990 590 1050 605
rect 990 570 1010 590
rect 1030 570 1050 590
rect 770 550 830 565
rect 880 550 940 565
rect 990 550 1050 570
rect 1100 590 1160 605
rect 1100 570 1120 590
rect 1140 570 1160 590
rect 1100 550 1160 570
rect 1210 590 1270 605
rect 1210 570 1230 590
rect 1250 570 1270 590
rect 1210 550 1270 570
rect 1320 590 1380 605
rect 1320 570 1340 590
rect 1360 570 1380 590
rect 1320 550 1380 570
rect 0 190 60 400
rect 0 170 20 190
rect 40 170 60 190
rect 0 150 60 170
rect 110 270 170 400
rect 220 385 280 400
rect 110 250 130 270
rect 150 250 170 270
rect 110 150 170 250
rect 220 270 280 280
rect 220 250 240 270
rect 260 250 280 270
rect 220 150 280 250
rect 330 270 390 400
rect 330 250 350 270
rect 370 250 390 270
rect 330 150 390 250
rect 440 240 500 400
rect 550 240 610 400
rect 660 385 720 400
rect 770 205 830 400
rect 880 205 940 400
rect 990 385 1050 400
rect 1100 385 1160 400
rect 1210 385 1270 400
rect 1320 385 1380 400
rect 440 190 610 205
rect 440 170 515 190
rect 535 170 610 190
rect 440 160 610 170
rect 440 150 500 160
rect 550 150 610 160
rect 660 190 720 205
rect 660 170 680 190
rect 700 170 720 190
rect 660 150 720 170
rect 770 190 940 205
rect 770 170 900 190
rect 920 170 940 190
rect 770 160 940 170
rect 770 150 830 160
rect 880 150 940 160
rect 990 190 1050 205
rect 990 170 1010 190
rect 1030 170 1050 190
rect 990 150 1050 170
rect 1100 190 1160 205
rect 1100 170 1120 190
rect 1140 170 1160 190
rect 1100 150 1160 170
rect 1210 190 1270 205
rect 1210 170 1230 190
rect 1250 170 1270 190
rect 1210 150 1270 170
rect 1320 190 1380 205
rect 1320 170 1340 190
rect 1360 170 1380 190
rect 1320 150 1380 170
rect 0 -15 60 0
rect 110 -15 170 0
rect 220 -15 280 0
rect 330 -15 390 0
rect 440 -15 500 0
rect 550 -15 610 0
rect 660 -15 720 0
rect 770 -15 830 0
rect 880 -15 940 0
rect 990 -15 1050 0
rect 1100 -15 1160 0
rect 1210 -15 1270 0
rect 1320 -15 1380 0
<< polycont >>
rect 240 570 260 590
rect 680 570 700 590
rect 1010 570 1030 590
rect 1120 570 1140 590
rect 1230 570 1250 590
rect 1340 570 1360 590
rect 20 170 40 190
rect 130 250 150 270
rect 240 250 260 270
rect 350 250 370 270
rect 515 170 535 190
rect 680 170 700 190
rect 900 170 920 190
rect 1010 170 1030 190
rect 1120 170 1140 190
rect 1230 170 1250 190
rect 1340 170 1360 190
<< locali >>
rect -95 535 -5 545
rect -95 415 -85 535
rect -65 415 -35 535
rect -15 415 -5 535
rect -95 200 -5 415
rect 65 535 105 715
rect 230 590 270 600
rect 230 570 240 590
rect 260 570 270 590
rect 230 560 270 570
rect 290 545 320 715
rect 670 590 710 720
rect 670 570 680 590
rect 700 570 710 590
rect 670 560 710 570
rect 730 545 760 720
rect 65 415 75 535
rect 95 415 105 535
rect 65 405 105 415
rect 175 535 215 545
rect 175 415 185 535
rect 205 415 215 535
rect 175 280 215 415
rect 285 535 325 545
rect 285 415 295 535
rect 315 415 325 535
rect 285 405 325 415
rect 395 535 435 545
rect 395 415 405 535
rect 425 415 435 535
rect 395 405 435 415
rect 505 535 545 545
rect 505 415 515 535
rect 535 415 545 535
rect 505 405 545 415
rect 615 535 655 545
rect 615 415 625 535
rect 645 415 655 535
rect 615 405 655 415
rect 725 535 765 545
rect 725 415 735 535
rect 755 415 765 535
rect 725 405 765 415
rect 120 270 270 280
rect 120 250 130 270
rect 150 250 185 270
rect 205 250 240 270
rect 260 250 270 270
rect 120 240 270 250
rect 340 270 380 280
rect 340 250 350 270
rect 370 250 380 270
rect 340 240 380 250
rect -95 190 50 200
rect -95 170 20 190
rect 40 170 50 190
rect 400 185 430 405
rect 450 270 490 280
rect 450 250 460 270
rect 480 250 490 270
rect 450 240 490 250
rect 510 205 540 405
rect 560 270 600 280
rect 560 250 570 270
rect 590 250 600 270
rect 560 240 600 250
rect -95 160 50 170
rect 175 165 430 185
rect -95 135 -5 160
rect -95 15 -85 135
rect -65 15 -35 135
rect -15 15 -5 135
rect -95 5 -5 15
rect 65 135 105 145
rect 65 15 75 135
rect 95 15 105 135
rect 65 -65 105 15
rect 175 135 215 165
rect 395 145 430 165
rect 505 190 545 205
rect 505 170 515 190
rect 535 170 545 190
rect 175 15 185 135
rect 205 15 215 135
rect 175 5 215 15
rect 285 135 325 145
rect 285 15 295 135
rect 315 15 325 135
rect 65 -85 75 -65
rect 95 -85 105 -65
rect 65 -95 105 -85
rect 285 -65 325 15
rect 395 135 435 145
rect 395 15 405 135
rect 425 15 435 135
rect 395 5 435 15
rect 505 135 545 170
rect 620 145 650 405
rect 670 195 710 200
rect 785 195 815 720
rect 670 190 815 195
rect 670 170 680 190
rect 700 170 815 190
rect 670 165 815 170
rect 670 160 710 165
rect 840 145 870 720
rect 1000 590 1040 600
rect 1000 570 1010 590
rect 1030 570 1040 590
rect 1000 560 1040 570
rect 1110 590 1150 600
rect 1110 570 1120 590
rect 1140 570 1150 590
rect 1110 560 1150 570
rect 1220 590 1260 600
rect 1220 570 1230 590
rect 1250 570 1260 590
rect 1220 560 1260 570
rect 1330 590 1370 600
rect 1330 570 1340 590
rect 1360 570 1370 590
rect 1330 560 1370 570
rect 945 535 985 545
rect 945 415 955 535
rect 975 415 985 535
rect 945 405 985 415
rect 1055 535 1095 545
rect 1055 415 1065 535
rect 1085 415 1095 535
rect 1055 405 1095 415
rect 1165 535 1205 545
rect 1165 415 1175 535
rect 1195 415 1205 535
rect 1165 405 1205 415
rect 1275 535 1315 545
rect 1275 415 1285 535
rect 1305 415 1315 535
rect 1275 405 1315 415
rect 1385 535 1480 545
rect 1385 415 1395 535
rect 1415 415 1445 535
rect 1465 415 1480 535
rect 1385 405 1480 415
rect 890 190 930 200
rect 890 170 900 190
rect 920 170 930 190
rect 890 160 930 170
rect 1000 190 1040 200
rect 1000 170 1010 190
rect 1030 170 1040 190
rect 1000 160 1040 170
rect 1110 190 1150 200
rect 1110 170 1120 190
rect 1140 170 1150 190
rect 1110 160 1150 170
rect 1220 190 1260 200
rect 1220 170 1230 190
rect 1250 170 1260 190
rect 1220 160 1260 170
rect 1330 190 1370 200
rect 1330 170 1340 190
rect 1360 170 1370 190
rect 1330 160 1370 170
rect 505 15 515 135
rect 535 15 545 135
rect 505 5 545 15
rect 615 135 655 145
rect 615 15 625 135
rect 645 15 655 135
rect 615 5 655 15
rect 725 135 870 145
rect 725 15 735 135
rect 755 115 870 135
rect 945 135 985 145
rect 755 15 765 115
rect 725 5 765 15
rect 945 15 955 135
rect 975 15 985 135
rect 945 5 985 15
rect 1055 135 1095 145
rect 1055 15 1065 135
rect 1085 15 1095 135
rect 1055 5 1095 15
rect 1165 135 1205 145
rect 1165 15 1175 135
rect 1195 15 1205 135
rect 1165 5 1205 15
rect 1275 135 1315 145
rect 1275 15 1285 135
rect 1305 15 1315 135
rect 1275 5 1315 15
rect 1385 135 1480 145
rect 1385 15 1395 135
rect 1415 15 1445 135
rect 1465 15 1480 135
rect 1385 5 1480 15
rect 285 -85 295 -65
rect 315 -85 325 -65
rect 285 -95 325 -85
<< viali >>
rect -85 415 -65 535
rect -35 415 -15 535
rect 240 570 260 590
rect 515 415 535 535
rect 130 250 150 270
rect 185 250 205 270
rect 240 250 260 270
rect 350 250 370 270
rect 460 250 480 270
rect 570 250 590 270
rect -85 15 -65 135
rect -35 15 -15 135
rect 75 -85 95 -65
rect 900 170 920 190
rect 515 15 535 135
rect 295 -85 315 -65
<< metal1 >>
rect 230 590 270 600
rect 230 570 240 590
rect 260 570 270 590
rect 230 545 270 570
rect -100 535 1480 545
rect -100 415 -85 535
rect -65 415 -35 535
rect -15 415 515 535
rect 535 415 1480 535
rect -100 405 1480 415
rect -100 270 1485 280
rect -100 250 130 270
rect 150 250 185 270
rect 205 250 240 270
rect 260 250 350 270
rect 370 250 460 270
rect 480 250 570 270
rect 590 250 1485 270
rect -100 240 1485 250
rect 890 190 930 200
rect 890 170 900 190
rect 920 170 930 190
rect 890 145 930 170
rect -100 135 1480 145
rect -100 15 -85 135
rect -65 15 -35 135
rect -15 15 515 135
rect 535 15 1480 135
rect -100 5 1480 15
rect -100 -65 1480 -55
rect -100 -85 75 -65
rect 95 -85 295 -65
rect 315 -85 1480 -65
rect -100 -95 1480 -85
<< end >>
