magic
tech sky130A
timestamp 1620794316
<< nwell >>
rect -90 205 450 345
<< nmos >>
rect 95 70 110 170
rect 160 70 175 170
<< pmos >>
rect 30 225 45 325
rect 95 225 110 325
rect 250 225 265 325
rect 315 225 330 325
<< ndiff >>
rect 45 155 95 170
rect 45 85 60 155
rect 80 85 95 155
rect 45 70 95 85
rect 110 70 160 170
rect 175 155 230 170
rect 175 85 195 155
rect 215 85 230 155
rect 175 70 230 85
<< pdiff >>
rect -20 310 30 325
rect -20 240 -5 310
rect 15 240 30 310
rect -20 225 30 240
rect 45 310 95 325
rect 45 240 60 310
rect 80 240 95 310
rect 45 225 95 240
rect 110 310 160 325
rect 110 240 125 310
rect 145 240 160 310
rect 110 225 160 240
rect 200 310 250 325
rect 200 240 215 310
rect 235 240 250 310
rect 200 225 250 240
rect 265 310 315 325
rect 265 240 280 310
rect 300 240 315 310
rect 265 225 315 240
rect 330 310 380 325
rect 330 240 345 310
rect 365 240 380 310
rect 330 225 380 240
<< ndiffc >>
rect 60 85 80 155
rect 195 85 215 155
<< pdiffc >>
rect -5 240 15 310
rect 60 240 80 310
rect 125 240 145 310
rect 215 240 235 310
rect 280 240 300 310
rect 345 240 365 310
<< psubdiff >>
rect -5 155 45 170
rect -5 85 10 155
rect 30 85 45 155
rect -5 70 45 85
<< nsubdiff >>
rect -70 310 -20 325
rect -70 240 -55 310
rect -35 240 -20 310
rect -70 225 -20 240
rect 380 310 430 325
rect 380 240 395 310
rect 415 240 430 310
rect 380 225 430 240
<< psubdiffcont >>
rect 10 85 30 155
<< nsubdiffcont >>
rect -55 240 -35 310
rect 395 240 415 310
<< poly >>
rect 30 325 45 340
rect 95 325 110 340
rect 250 325 265 340
rect 315 325 330 340
rect 30 210 45 225
rect 95 210 110 225
rect 250 210 265 225
rect 315 210 330 225
rect 30 195 110 210
rect 95 170 110 195
rect 160 195 330 210
rect 160 170 175 195
rect 95 55 110 70
rect 160 55 175 70
rect 70 45 110 55
rect 70 25 80 45
rect 100 25 110 45
rect 70 15 110 25
rect 135 45 175 55
rect 135 25 145 45
rect 165 25 175 45
rect 135 15 175 25
<< polycont >>
rect 80 25 100 45
rect 145 25 165 45
<< locali >>
rect -65 310 25 320
rect -65 240 -55 310
rect -35 240 -5 310
rect 15 240 25 310
rect -65 230 25 240
rect 50 310 90 320
rect 50 240 60 310
rect 80 240 90 310
rect 50 230 90 240
rect 115 310 155 320
rect 115 240 125 310
rect 145 240 155 310
rect 115 230 155 240
rect 205 310 245 320
rect 205 240 215 310
rect 235 240 245 310
rect 205 230 245 240
rect 270 310 310 320
rect 270 240 280 310
rect 300 240 310 310
rect 270 230 310 240
rect 335 310 425 320
rect 335 240 345 310
rect 365 240 395 310
rect 415 240 425 310
rect 335 230 425 240
rect 70 205 90 230
rect 270 205 290 230
rect 70 185 290 205
rect 205 165 225 185
rect 0 155 90 165
rect 0 85 10 155
rect 30 85 60 155
rect 80 85 90 155
rect 0 75 90 85
rect 185 155 225 165
rect 185 85 195 155
rect 215 85 225 155
rect 185 75 225 85
rect 205 55 225 75
rect 70 45 110 55
rect 70 25 80 45
rect 100 25 110 45
rect 70 15 110 25
rect 135 45 175 55
rect 135 25 145 45
rect 165 25 175 45
rect 205 35 385 55
rect 135 15 175 25
rect 80 0 100 15
rect 145 0 165 15
<< viali >>
rect -55 240 -35 310
rect -5 240 15 310
rect 125 240 145 310
rect 215 240 235 310
rect 345 240 365 310
rect 395 240 415 310
rect 10 85 30 155
rect 60 85 80 155
<< metal1 >>
rect -90 310 450 320
rect -90 240 -55 310
rect -35 240 -5 310
rect 15 240 125 310
rect 145 240 215 310
rect 235 240 345 310
rect 365 240 395 310
rect 415 240 450 310
rect -90 230 450 240
rect -25 155 250 165
rect -25 85 10 155
rect 30 85 60 155
rect 80 85 250 155
rect -25 75 250 85
<< labels >>
rlabel locali 90 0 90 0 5 A
port 1 s
rlabel locali 155 0 155 0 5 B
port 2 s
rlabel locali 385 45 385 45 5 Y
port 3 s
rlabel metal1 -25 120 -25 120 7 VN
port 4 w
rlabel metal1 -90 275 -90 275 7 VP
port 5 w
rlabel ndiff 135 115 135 115 5 net1
<< end >>
