magic
tech sky130A
timestamp 1620673804
<< xpolycontact >>
rect 0 1095 35 1315
rect 0 0 35 220
rect 160 1095 195 1315
rect 160 0 195 220
rect 320 1095 355 1315
rect 320 0 355 220
rect 480 1095 515 1315
rect 480 0 515 220
rect 640 1095 675 1315
rect 640 0 675 220
<< xpolyres >>
rect 0 220 35 1095
rect 160 220 195 1095
rect 320 220 355 1095
rect 480 220 515 1095
rect 640 220 675 1095
<< locali >>
rect 35 1095 160 1315
rect 355 1095 480 1315
rect 195 0 320 220
rect 515 0 640 220
<< end >>
