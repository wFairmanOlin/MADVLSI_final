magic
tech sky130A
timestamp 1620822988
<< nwell >>
rect -120 1150 3030 1670
<< nmos >>
rect 0 400 60 550
rect 110 400 170 550
rect 220 400 280 550
rect 330 400 390 550
rect 440 400 500 550
rect 550 400 610 550
rect 660 400 720 550
rect 770 400 830 550
rect 880 400 940 550
rect 990 400 1050 550
rect 1100 400 1160 550
rect 1210 400 1270 550
rect 1320 400 1380 550
rect 1530 400 1590 550
rect 1640 400 1700 550
rect 1750 400 1810 550
rect 1860 400 1920 550
rect 1970 400 2030 550
rect 2080 400 2140 550
rect 2190 400 2250 550
rect 2300 400 2360 550
rect 2410 400 2470 550
rect 2520 400 2580 550
rect 2630 400 2690 550
rect 2740 400 2800 550
rect 2850 400 2910 550
rect 0 80 60 230
rect 110 80 170 230
rect 220 80 280 230
rect 330 80 390 230
rect 440 80 500 230
rect 550 80 610 230
rect 660 80 720 230
rect 770 80 830 230
rect 880 80 940 230
rect 990 80 1050 230
rect 1100 80 1160 230
rect 1210 80 1270 230
rect 1320 80 1380 230
rect 1530 80 1590 230
rect 1640 80 1700 230
rect 1750 80 1810 230
rect 1860 80 1920 230
rect 1970 80 2030 230
rect 2080 80 2140 230
rect 2190 80 2250 230
rect 2300 80 2360 230
rect 2410 80 2470 230
rect 2520 80 2580 230
rect 2630 80 2690 230
rect 2740 80 2800 230
rect 2850 80 2910 230
<< pmos >>
rect 0 1500 60 1650
rect 110 1500 170 1650
rect 220 1500 280 1650
rect 330 1500 390 1650
rect 440 1500 500 1650
rect 550 1500 610 1650
rect 660 1500 720 1650
rect 770 1500 830 1650
rect 880 1500 940 1650
rect 990 1500 1050 1650
rect 1100 1500 1160 1650
rect 1210 1500 1270 1650
rect 1320 1500 1380 1650
rect 1530 1500 1590 1650
rect 1640 1500 1700 1650
rect 1750 1500 1810 1650
rect 1860 1500 1920 1650
rect 1970 1500 2030 1650
rect 2080 1500 2140 1650
rect 2190 1500 2250 1650
rect 2300 1500 2360 1650
rect 2410 1500 2470 1650
rect 2520 1500 2580 1650
rect 2630 1500 2690 1650
rect 2740 1500 2800 1650
rect 2850 1500 2910 1650
rect 0 1170 60 1320
rect 110 1170 170 1320
rect 220 1170 280 1320
rect 330 1170 390 1320
rect 440 1170 500 1320
rect 550 1170 610 1320
rect 660 1170 720 1320
rect 770 1170 830 1320
rect 880 1170 940 1320
rect 990 1170 1050 1320
rect 1100 1170 1160 1320
rect 1210 1170 1270 1320
rect 1320 1170 1380 1320
rect 1530 1170 1590 1320
rect 1640 1170 1700 1320
rect 1750 1170 1810 1320
rect 1860 1170 1920 1320
rect 1970 1170 2030 1320
rect 2080 1170 2140 1320
rect 2190 1170 2250 1320
rect 2300 1170 2360 1320
rect 2410 1170 2470 1320
rect 2520 1170 2580 1320
rect 2630 1170 2690 1320
rect 2740 1170 2800 1320
rect 2850 1170 2910 1320
<< ndiff >>
rect -50 535 0 550
rect -50 415 -35 535
rect -15 415 0 535
rect -50 400 0 415
rect 60 535 110 550
rect 60 415 75 535
rect 95 415 110 535
rect 60 400 110 415
rect 170 535 220 550
rect 170 415 185 535
rect 205 415 220 535
rect 170 400 220 415
rect 280 535 330 550
rect 280 415 295 535
rect 315 415 330 535
rect 280 400 330 415
rect 390 535 440 550
rect 390 415 405 535
rect 425 415 440 535
rect 390 400 440 415
rect 500 535 550 550
rect 500 415 515 535
rect 535 415 550 535
rect 500 400 550 415
rect 610 535 660 550
rect 610 415 625 535
rect 645 415 660 535
rect 610 400 660 415
rect 720 535 770 550
rect 720 415 735 535
rect 755 415 770 535
rect 720 400 770 415
rect 830 400 880 550
rect 940 535 990 550
rect 940 415 955 535
rect 975 415 990 535
rect 940 400 990 415
rect 1050 535 1100 550
rect 1050 415 1065 535
rect 1085 415 1100 535
rect 1050 400 1100 415
rect 1160 535 1210 550
rect 1160 415 1175 535
rect 1195 415 1210 535
rect 1160 400 1210 415
rect 1270 535 1320 550
rect 1270 415 1285 535
rect 1305 415 1320 535
rect 1270 400 1320 415
rect 1380 535 1430 550
rect 1480 535 1530 550
rect 1380 415 1395 535
rect 1415 415 1430 535
rect 1480 415 1495 535
rect 1515 415 1530 535
rect 1380 400 1430 415
rect 1480 400 1530 415
rect 1590 535 1640 550
rect 1590 415 1605 535
rect 1625 415 1640 535
rect 1590 400 1640 415
rect 1700 535 1750 550
rect 1700 415 1715 535
rect 1735 415 1750 535
rect 1700 400 1750 415
rect 1810 535 1860 550
rect 1810 415 1825 535
rect 1845 415 1860 535
rect 1810 400 1860 415
rect 1920 535 1970 550
rect 1920 415 1935 535
rect 1955 415 1970 535
rect 1920 400 1970 415
rect 2030 400 2080 550
rect 2140 535 2190 550
rect 2140 415 2155 535
rect 2175 415 2190 535
rect 2140 400 2190 415
rect 2250 535 2300 550
rect 2250 415 2265 535
rect 2285 415 2300 535
rect 2250 400 2300 415
rect 2360 535 2410 550
rect 2360 415 2375 535
rect 2395 415 2410 535
rect 2360 400 2410 415
rect 2470 535 2520 550
rect 2470 415 2485 535
rect 2505 415 2520 535
rect 2470 400 2520 415
rect 2580 535 2630 550
rect 2580 415 2595 535
rect 2615 415 2630 535
rect 2580 400 2630 415
rect 2690 535 2740 550
rect 2690 415 2705 535
rect 2725 415 2740 535
rect 2690 400 2740 415
rect 2800 535 2850 550
rect 2800 415 2815 535
rect 2835 415 2850 535
rect 2800 400 2850 415
rect 2910 535 2960 550
rect 2910 415 2925 535
rect 2945 415 2960 535
rect 2910 400 2960 415
rect -50 215 0 230
rect -50 95 -35 215
rect -15 95 0 215
rect -50 80 0 95
rect 60 215 110 230
rect 60 95 75 215
rect 95 95 110 215
rect 60 80 110 95
rect 170 215 220 230
rect 170 95 185 215
rect 205 95 220 215
rect 170 80 220 95
rect 280 215 330 230
rect 280 95 295 215
rect 315 95 330 215
rect 280 80 330 95
rect 390 215 440 230
rect 390 95 405 215
rect 425 95 440 215
rect 390 80 440 95
rect 500 215 550 230
rect 500 95 515 215
rect 535 95 550 215
rect 500 80 550 95
rect 610 215 660 230
rect 610 95 625 215
rect 645 95 660 215
rect 610 80 660 95
rect 720 215 770 230
rect 720 95 735 215
rect 755 95 770 215
rect 720 80 770 95
rect 830 80 880 230
rect 940 215 990 230
rect 940 95 955 215
rect 975 95 990 215
rect 940 80 990 95
rect 1050 215 1100 230
rect 1050 95 1065 215
rect 1085 95 1100 215
rect 1050 80 1100 95
rect 1160 215 1210 230
rect 1160 95 1175 215
rect 1195 95 1210 215
rect 1160 80 1210 95
rect 1270 215 1320 230
rect 1270 95 1285 215
rect 1305 95 1320 215
rect 1270 80 1320 95
rect 1380 215 1430 230
rect 1480 215 1530 230
rect 1380 95 1395 215
rect 1415 95 1430 215
rect 1480 95 1495 215
rect 1515 95 1530 215
rect 1380 80 1430 95
rect 1480 80 1530 95
rect 1590 215 1640 230
rect 1590 95 1605 215
rect 1625 95 1640 215
rect 1590 80 1640 95
rect 1700 215 1750 230
rect 1700 95 1715 215
rect 1735 95 1750 215
rect 1700 80 1750 95
rect 1810 215 1860 230
rect 1810 95 1825 215
rect 1845 95 1860 215
rect 1810 80 1860 95
rect 1920 215 1970 230
rect 1920 95 1935 215
rect 1955 95 1970 215
rect 1920 80 1970 95
rect 2030 80 2080 230
rect 2140 215 2190 230
rect 2140 95 2155 215
rect 2175 95 2190 215
rect 2140 80 2190 95
rect 2250 215 2300 230
rect 2250 95 2265 215
rect 2285 95 2300 215
rect 2250 80 2300 95
rect 2360 215 2410 230
rect 2360 95 2375 215
rect 2395 95 2410 215
rect 2360 80 2410 95
rect 2470 215 2520 230
rect 2470 95 2485 215
rect 2505 95 2520 215
rect 2470 80 2520 95
rect 2580 215 2630 230
rect 2580 95 2595 215
rect 2615 95 2630 215
rect 2580 80 2630 95
rect 2690 215 2740 230
rect 2690 95 2705 215
rect 2725 95 2740 215
rect 2690 80 2740 95
rect 2800 215 2850 230
rect 2800 95 2815 215
rect 2835 95 2850 215
rect 2800 80 2850 95
rect 2910 215 2960 230
rect 2910 95 2925 215
rect 2945 95 2960 215
rect 2910 80 2960 95
<< pdiff >>
rect -50 1635 0 1650
rect -50 1515 -35 1635
rect -15 1515 0 1635
rect -50 1500 0 1515
rect 60 1635 110 1650
rect 60 1515 75 1635
rect 95 1515 110 1635
rect 60 1500 110 1515
rect 170 1635 220 1650
rect 170 1515 185 1635
rect 205 1515 220 1635
rect 170 1500 220 1515
rect 280 1635 330 1650
rect 280 1515 295 1635
rect 315 1515 330 1635
rect 280 1500 330 1515
rect 390 1635 440 1650
rect 390 1515 405 1635
rect 425 1515 440 1635
rect 390 1500 440 1515
rect 500 1635 550 1650
rect 500 1515 515 1635
rect 535 1515 550 1635
rect 500 1500 550 1515
rect 610 1635 660 1650
rect 610 1515 625 1635
rect 645 1515 660 1635
rect 610 1500 660 1515
rect 720 1635 770 1650
rect 720 1515 735 1635
rect 755 1515 770 1635
rect 720 1500 770 1515
rect 830 1500 880 1650
rect 940 1635 990 1650
rect 940 1515 955 1635
rect 975 1515 990 1635
rect 940 1500 990 1515
rect 1050 1635 1100 1650
rect 1050 1515 1065 1635
rect 1085 1515 1100 1635
rect 1050 1500 1100 1515
rect 1160 1635 1210 1650
rect 1160 1515 1175 1635
rect 1195 1515 1210 1635
rect 1160 1500 1210 1515
rect 1270 1635 1320 1650
rect 1270 1515 1285 1635
rect 1305 1515 1320 1635
rect 1270 1500 1320 1515
rect 1380 1635 1430 1650
rect 1480 1635 1530 1650
rect 1380 1515 1395 1635
rect 1415 1515 1430 1635
rect 1480 1515 1495 1635
rect 1515 1515 1530 1635
rect 1380 1500 1430 1515
rect 1480 1500 1530 1515
rect 1590 1635 1640 1650
rect 1590 1515 1605 1635
rect 1625 1515 1640 1635
rect 1590 1500 1640 1515
rect 1700 1635 1750 1650
rect 1700 1515 1715 1635
rect 1735 1515 1750 1635
rect 1700 1500 1750 1515
rect 1810 1635 1860 1650
rect 1810 1515 1825 1635
rect 1845 1515 1860 1635
rect 1810 1500 1860 1515
rect 1920 1635 1970 1650
rect 1920 1515 1935 1635
rect 1955 1515 1970 1635
rect 1920 1500 1970 1515
rect 2030 1500 2080 1650
rect 2140 1635 2190 1650
rect 2140 1515 2155 1635
rect 2175 1515 2190 1635
rect 2140 1500 2190 1515
rect 2250 1635 2300 1650
rect 2250 1515 2265 1635
rect 2285 1515 2300 1635
rect 2250 1500 2300 1515
rect 2360 1635 2410 1650
rect 2360 1515 2375 1635
rect 2395 1515 2410 1635
rect 2360 1500 2410 1515
rect 2470 1635 2520 1650
rect 2470 1515 2485 1635
rect 2505 1515 2520 1635
rect 2470 1500 2520 1515
rect 2580 1635 2630 1650
rect 2580 1515 2595 1635
rect 2615 1515 2630 1635
rect 2580 1500 2630 1515
rect 2690 1635 2740 1650
rect 2690 1515 2705 1635
rect 2725 1515 2740 1635
rect 2690 1500 2740 1515
rect 2800 1635 2850 1650
rect 2800 1515 2815 1635
rect 2835 1515 2850 1635
rect 2800 1500 2850 1515
rect 2910 1635 2960 1650
rect 2910 1515 2925 1635
rect 2945 1515 2960 1635
rect 2910 1500 2960 1515
rect -50 1305 0 1320
rect -50 1185 -35 1305
rect -15 1185 0 1305
rect -50 1170 0 1185
rect 60 1305 110 1320
rect 60 1185 75 1305
rect 95 1185 110 1305
rect 60 1170 110 1185
rect 170 1305 220 1320
rect 170 1185 185 1305
rect 205 1185 220 1305
rect 170 1170 220 1185
rect 280 1305 330 1320
rect 280 1185 295 1305
rect 315 1185 330 1305
rect 280 1170 330 1185
rect 390 1305 440 1320
rect 390 1185 405 1305
rect 425 1185 440 1305
rect 390 1170 440 1185
rect 500 1305 550 1320
rect 500 1185 515 1305
rect 535 1185 550 1305
rect 500 1170 550 1185
rect 610 1305 660 1320
rect 610 1185 625 1305
rect 645 1185 660 1305
rect 610 1170 660 1185
rect 720 1305 770 1320
rect 720 1185 735 1305
rect 755 1185 770 1305
rect 720 1170 770 1185
rect 830 1170 880 1320
rect 940 1305 990 1320
rect 940 1185 955 1305
rect 975 1185 990 1305
rect 940 1170 990 1185
rect 1050 1305 1100 1320
rect 1050 1185 1065 1305
rect 1085 1185 1100 1305
rect 1050 1170 1100 1185
rect 1160 1305 1210 1320
rect 1160 1185 1175 1305
rect 1195 1185 1210 1305
rect 1160 1170 1210 1185
rect 1270 1305 1320 1320
rect 1270 1185 1285 1305
rect 1305 1185 1320 1305
rect 1270 1170 1320 1185
rect 1380 1305 1430 1320
rect 1480 1305 1530 1320
rect 1380 1185 1395 1305
rect 1415 1185 1430 1305
rect 1480 1185 1495 1305
rect 1515 1185 1530 1305
rect 1380 1170 1430 1185
rect 1480 1170 1530 1185
rect 1590 1305 1640 1320
rect 1590 1185 1605 1305
rect 1625 1185 1640 1305
rect 1590 1170 1640 1185
rect 1700 1305 1750 1320
rect 1700 1185 1715 1305
rect 1735 1185 1750 1305
rect 1700 1170 1750 1185
rect 1810 1305 1860 1320
rect 1810 1185 1825 1305
rect 1845 1185 1860 1305
rect 1810 1170 1860 1185
rect 1920 1305 1970 1320
rect 1920 1185 1935 1305
rect 1955 1185 1970 1305
rect 1920 1170 1970 1185
rect 2030 1170 2080 1320
rect 2140 1305 2190 1320
rect 2140 1185 2155 1305
rect 2175 1185 2190 1305
rect 2140 1170 2190 1185
rect 2250 1305 2300 1320
rect 2250 1185 2265 1305
rect 2285 1185 2300 1305
rect 2250 1170 2300 1185
rect 2360 1305 2410 1320
rect 2360 1185 2375 1305
rect 2395 1185 2410 1305
rect 2360 1170 2410 1185
rect 2470 1305 2520 1320
rect 2470 1185 2485 1305
rect 2505 1185 2520 1305
rect 2470 1170 2520 1185
rect 2580 1305 2630 1320
rect 2580 1185 2595 1305
rect 2615 1185 2630 1305
rect 2580 1170 2630 1185
rect 2690 1305 2740 1320
rect 2690 1185 2705 1305
rect 2725 1185 2740 1305
rect 2690 1170 2740 1185
rect 2800 1305 2850 1320
rect 2800 1185 2815 1305
rect 2835 1185 2850 1305
rect 2800 1170 2850 1185
rect 2910 1305 2960 1320
rect 2910 1185 2925 1305
rect 2945 1185 2960 1305
rect 2910 1170 2960 1185
<< ndiffc >>
rect -35 415 -15 535
rect 75 415 95 535
rect 185 415 205 535
rect 295 415 315 535
rect 405 415 425 535
rect 515 415 535 535
rect 625 415 645 535
rect 735 415 755 535
rect 955 415 975 535
rect 1065 415 1085 535
rect 1175 415 1195 535
rect 1285 415 1305 535
rect 1395 415 1415 535
rect 1495 415 1515 535
rect 1605 415 1625 535
rect 1715 415 1735 535
rect 1825 415 1845 535
rect 1935 415 1955 535
rect 2155 415 2175 535
rect 2265 415 2285 535
rect 2375 415 2395 535
rect 2485 415 2505 535
rect 2595 415 2615 535
rect 2705 415 2725 535
rect 2815 415 2835 535
rect 2925 415 2945 535
rect -35 95 -15 215
rect 75 95 95 215
rect 185 95 205 215
rect 295 95 315 215
rect 405 95 425 215
rect 515 95 535 215
rect 625 95 645 215
rect 735 95 755 215
rect 955 95 975 215
rect 1065 95 1085 215
rect 1175 95 1195 215
rect 1285 95 1305 215
rect 1395 95 1415 215
rect 1495 95 1515 215
rect 1605 95 1625 215
rect 1715 95 1735 215
rect 1825 95 1845 215
rect 1935 95 1955 215
rect 2155 95 2175 215
rect 2265 95 2285 215
rect 2375 95 2395 215
rect 2485 95 2505 215
rect 2595 95 2615 215
rect 2705 95 2725 215
rect 2815 95 2835 215
rect 2925 95 2945 215
<< pdiffc >>
rect -35 1515 -15 1635
rect 75 1515 95 1635
rect 185 1515 205 1635
rect 295 1515 315 1635
rect 405 1515 425 1635
rect 515 1515 535 1635
rect 625 1515 645 1635
rect 735 1515 755 1635
rect 955 1515 975 1635
rect 1065 1515 1085 1635
rect 1175 1515 1195 1635
rect 1285 1515 1305 1635
rect 1395 1515 1415 1635
rect 1495 1515 1515 1635
rect 1605 1515 1625 1635
rect 1715 1515 1735 1635
rect 1825 1515 1845 1635
rect 1935 1515 1955 1635
rect 2155 1515 2175 1635
rect 2265 1515 2285 1635
rect 2375 1515 2395 1635
rect 2485 1515 2505 1635
rect 2595 1515 2615 1635
rect 2705 1515 2725 1635
rect 2815 1515 2835 1635
rect 2925 1515 2945 1635
rect -35 1185 -15 1305
rect 75 1185 95 1305
rect 185 1185 205 1305
rect 295 1185 315 1305
rect 405 1185 425 1305
rect 515 1185 535 1305
rect 625 1185 645 1305
rect 735 1185 755 1305
rect 955 1185 975 1305
rect 1065 1185 1085 1305
rect 1175 1185 1195 1305
rect 1285 1185 1305 1305
rect 1395 1185 1415 1305
rect 1495 1185 1515 1305
rect 1605 1185 1625 1305
rect 1715 1185 1735 1305
rect 1825 1185 1845 1305
rect 1935 1185 1955 1305
rect 2155 1185 2175 1305
rect 2265 1185 2285 1305
rect 2375 1185 2395 1305
rect 2485 1185 2505 1305
rect 2595 1185 2615 1305
rect 2705 1185 2725 1305
rect 2815 1185 2835 1305
rect 2925 1185 2945 1305
<< psubdiff >>
rect -100 535 -50 550
rect -100 415 -85 535
rect -65 415 -50 535
rect -100 400 -50 415
rect 1430 535 1480 550
rect 1430 415 1445 535
rect 1465 415 1480 535
rect 1430 400 1480 415
rect 2960 535 3010 550
rect 2960 415 2975 535
rect 2995 415 3010 535
rect 2960 400 3010 415
rect -100 215 -50 230
rect -100 95 -85 215
rect -65 95 -50 215
rect -100 80 -50 95
rect 1430 215 1480 230
rect 1430 95 1445 215
rect 1465 95 1480 215
rect 1430 80 1480 95
rect 2960 215 3010 230
rect 2960 95 2975 215
rect 2995 95 3010 215
rect 2960 80 3010 95
<< nsubdiff >>
rect -100 1635 -50 1650
rect -100 1515 -85 1635
rect -65 1515 -50 1635
rect -100 1500 -50 1515
rect 1430 1635 1480 1650
rect 1430 1515 1445 1635
rect 1465 1515 1480 1635
rect 1430 1500 1480 1515
rect 2960 1635 3010 1650
rect 2960 1515 2975 1635
rect 2995 1515 3010 1635
rect 2960 1500 3010 1515
rect -100 1305 -50 1320
rect -100 1185 -85 1305
rect -65 1185 -50 1305
rect -100 1170 -50 1185
rect 1430 1305 1480 1320
rect 1430 1185 1445 1305
rect 1465 1185 1480 1305
rect 1430 1170 1480 1185
rect 2960 1305 3010 1320
rect 2960 1185 2975 1305
rect 2995 1185 3010 1305
rect 2960 1170 3010 1185
<< psubdiffcont >>
rect -85 415 -65 535
rect 1445 415 1465 535
rect 2975 415 2995 535
rect -85 95 -65 215
rect 1445 95 1465 215
rect 2975 95 2995 215
<< nsubdiffcont >>
rect -85 1515 -65 1635
rect 1445 1515 1465 1635
rect 2975 1515 2995 1635
rect -85 1185 -65 1305
rect 1445 1185 1465 1305
rect 2975 1185 2995 1305
<< poly >>
rect 0 1650 60 1665
rect 110 1650 170 1665
rect 220 1650 280 1665
rect 330 1650 390 1665
rect 440 1650 500 1665
rect 550 1650 610 1665
rect 660 1650 720 1665
rect 770 1650 830 1665
rect 880 1650 940 1665
rect 990 1650 1050 1665
rect 1100 1650 1160 1665
rect 1210 1650 1270 1665
rect 1320 1650 1380 1665
rect 1530 1650 1590 1665
rect 1640 1650 1700 1665
rect 1750 1650 1810 1665
rect 1860 1650 1920 1665
rect 1970 1650 2030 1665
rect 2080 1650 2140 1665
rect 2190 1650 2250 1665
rect 2300 1650 2360 1665
rect 2410 1650 2470 1665
rect 2520 1650 2580 1665
rect 2630 1650 2690 1665
rect 2740 1650 2800 1665
rect 2850 1650 2910 1665
rect 0 1475 60 1500
rect 0 1455 20 1475
rect 40 1455 60 1475
rect 0 1320 60 1455
rect 110 1420 170 1500
rect 110 1400 130 1420
rect 150 1400 170 1420
rect 110 1320 170 1400
rect 220 1420 280 1500
rect 220 1400 240 1420
rect 260 1400 280 1420
rect 220 1390 280 1400
rect 330 1420 390 1500
rect 440 1485 500 1500
rect 550 1485 610 1500
rect 440 1475 610 1485
rect 440 1455 515 1475
rect 535 1455 610 1475
rect 440 1445 610 1455
rect 660 1475 720 1500
rect 660 1455 680 1475
rect 700 1455 720 1475
rect 660 1440 720 1455
rect 770 1485 830 1500
rect 880 1485 940 1500
rect 770 1475 940 1485
rect 770 1455 900 1475
rect 920 1455 940 1475
rect 770 1440 940 1455
rect 330 1400 350 1420
rect 370 1400 390 1420
rect 220 1320 280 1335
rect 330 1320 390 1400
rect 440 1365 500 1375
rect 440 1345 460 1365
rect 480 1345 500 1365
rect 440 1320 500 1345
rect 550 1365 610 1375
rect 550 1345 570 1365
rect 590 1345 610 1365
rect 550 1320 610 1345
rect 660 1320 720 1335
rect 770 1320 830 1440
rect 880 1320 940 1440
rect 990 1320 1050 1500
rect 1100 1420 1160 1500
rect 1100 1400 1120 1420
rect 1140 1400 1160 1420
rect 1100 1320 1160 1400
rect 1210 1320 1270 1500
rect 1320 1320 1380 1500
rect 1530 1320 1590 1500
rect 1640 1320 1700 1500
rect 1750 1420 1810 1500
rect 1750 1400 1770 1420
rect 1790 1400 1810 1420
rect 1750 1320 1810 1400
rect 1860 1320 1920 1500
rect 1970 1485 2030 1500
rect 2080 1485 2140 1500
rect 1970 1475 2140 1485
rect 1970 1455 1990 1475
rect 2010 1455 2140 1475
rect 1970 1440 2140 1455
rect 2190 1475 2250 1500
rect 2190 1455 2210 1475
rect 2230 1455 2250 1475
rect 2190 1440 2250 1455
rect 2300 1485 2360 1500
rect 2410 1485 2470 1500
rect 2300 1475 2470 1485
rect 2300 1455 2375 1475
rect 2395 1455 2470 1475
rect 2300 1445 2470 1455
rect 1970 1320 2030 1440
rect 2080 1320 2140 1440
rect 2520 1420 2580 1500
rect 2520 1400 2540 1420
rect 2560 1400 2580 1420
rect 2300 1365 2360 1375
rect 2300 1345 2320 1365
rect 2340 1345 2360 1365
rect 2190 1320 2250 1335
rect 2300 1320 2360 1345
rect 2410 1365 2470 1375
rect 2410 1345 2430 1365
rect 2450 1345 2470 1365
rect 2410 1320 2470 1345
rect 2520 1320 2580 1400
rect 2630 1420 2690 1500
rect 2630 1400 2650 1420
rect 2670 1400 2690 1420
rect 2630 1390 2690 1400
rect 2740 1420 2800 1500
rect 2740 1400 2760 1420
rect 2780 1400 2800 1420
rect 2630 1320 2690 1335
rect 2740 1320 2800 1400
rect 2850 1475 2910 1500
rect 2850 1455 2870 1475
rect 2890 1455 2910 1475
rect 2850 1320 2910 1455
rect 0 1150 60 1170
rect 110 1150 170 1170
rect 220 1145 280 1170
rect 330 1155 390 1170
rect 440 1155 500 1170
rect 550 1155 610 1170
rect 220 1125 240 1145
rect 260 1125 280 1145
rect 220 1110 280 1125
rect 660 1145 720 1170
rect 770 1150 830 1170
rect 880 1150 940 1170
rect 660 1125 680 1145
rect 700 1125 720 1145
rect 660 1110 720 1125
rect 990 1145 1050 1170
rect 1100 1150 1160 1170
rect 990 1125 1010 1145
rect 1030 1125 1050 1145
rect 990 1110 1050 1125
rect 1210 1145 1270 1170
rect 1210 1125 1230 1145
rect 1250 1125 1270 1145
rect 1210 1110 1270 1125
rect 1320 1145 1380 1170
rect 1320 1125 1340 1145
rect 1360 1125 1380 1145
rect 1320 1110 1380 1125
rect 1530 1145 1590 1170
rect 1530 1125 1550 1145
rect 1570 1125 1590 1145
rect 1530 1110 1590 1125
rect 1640 1145 1700 1170
rect 1750 1150 1810 1170
rect 1640 1125 1660 1145
rect 1680 1125 1700 1145
rect 1640 1110 1700 1125
rect 1860 1145 1920 1170
rect 1970 1150 2030 1170
rect 2080 1150 2140 1170
rect 1860 1125 1880 1145
rect 1900 1125 1920 1145
rect 1860 1110 1920 1125
rect 2190 1145 2250 1170
rect 2300 1155 2360 1170
rect 2410 1155 2470 1170
rect 2520 1155 2580 1170
rect 2190 1125 2210 1145
rect 2230 1125 2250 1145
rect 2190 1110 2250 1125
rect 2630 1145 2690 1170
rect 2740 1150 2800 1170
rect 2850 1150 2910 1170
rect 2630 1125 2650 1145
rect 2670 1125 2690 1145
rect 2630 1110 2690 1125
rect 220 590 280 605
rect 220 570 240 590
rect 260 570 280 590
rect 0 550 60 565
rect 110 550 170 565
rect 220 550 280 570
rect 660 590 720 605
rect 660 570 680 590
rect 700 570 720 590
rect 330 550 390 565
rect 440 550 500 565
rect 550 550 610 565
rect 660 550 720 570
rect 990 590 1050 605
rect 990 570 1010 590
rect 1030 570 1050 590
rect 770 550 830 565
rect 880 550 940 565
rect 990 550 1050 570
rect 1210 590 1270 605
rect 1210 570 1230 590
rect 1250 570 1270 590
rect 1100 550 1160 565
rect 1210 550 1270 570
rect 1320 590 1380 605
rect 1320 570 1340 590
rect 1360 570 1380 590
rect 1320 550 1380 570
rect 1530 590 1590 605
rect 1530 570 1550 590
rect 1570 570 1590 590
rect 1530 550 1590 570
rect 1640 590 1700 605
rect 1640 570 1660 590
rect 1680 570 1700 590
rect 1640 550 1700 570
rect 1860 590 1920 605
rect 1860 570 1880 590
rect 1900 570 1920 590
rect 1750 550 1810 565
rect 1860 550 1920 570
rect 2190 590 2250 605
rect 2190 570 2210 590
rect 2230 570 2250 590
rect 1970 550 2030 565
rect 2080 550 2140 565
rect 2190 550 2250 570
rect 2630 590 2690 605
rect 2630 570 2650 590
rect 2670 570 2690 590
rect 2300 550 2360 565
rect 2410 550 2470 565
rect 2520 550 2580 565
rect 2630 550 2690 570
rect 2740 550 2800 565
rect 2850 550 2910 565
rect 0 270 60 400
rect 0 250 20 270
rect 40 250 60 270
rect 0 230 60 250
rect 110 325 170 400
rect 220 385 280 400
rect 110 305 130 325
rect 150 305 170 325
rect 110 230 170 305
rect 220 325 280 335
rect 220 305 240 325
rect 260 305 280 325
rect 220 230 280 305
rect 330 325 390 400
rect 440 380 500 400
rect 440 360 460 380
rect 480 360 500 380
rect 440 350 500 360
rect 550 380 610 400
rect 660 385 720 400
rect 550 360 570 380
rect 590 360 610 380
rect 550 350 610 360
rect 330 305 350 325
rect 370 305 390 325
rect 330 230 390 305
rect 770 285 830 400
rect 880 285 940 400
rect 440 270 610 280
rect 440 250 515 270
rect 535 250 610 270
rect 440 240 610 250
rect 440 230 500 240
rect 550 230 610 240
rect 660 270 720 285
rect 660 250 680 270
rect 700 250 720 270
rect 660 230 720 250
rect 770 270 940 285
rect 770 250 900 270
rect 920 250 940 270
rect 770 240 940 250
rect 770 230 830 240
rect 880 230 940 240
rect 990 230 1050 400
rect 1100 325 1160 400
rect 1210 385 1270 400
rect 1100 305 1120 325
rect 1140 305 1160 325
rect 1100 230 1160 305
rect 1210 270 1270 285
rect 1210 250 1230 270
rect 1250 250 1270 270
rect 1210 230 1270 250
rect 1320 230 1380 400
rect 1530 230 1590 400
rect 1640 385 1700 400
rect 1750 325 1810 400
rect 1750 305 1770 325
rect 1790 305 1810 325
rect 1640 270 1700 285
rect 1640 250 1660 270
rect 1680 250 1700 270
rect 1640 230 1700 250
rect 1750 230 1810 305
rect 1860 230 1920 400
rect 1970 285 2030 400
rect 2080 285 2140 400
rect 2190 385 2250 400
rect 2300 380 2360 400
rect 2300 360 2320 380
rect 2340 360 2360 380
rect 2300 350 2360 360
rect 2410 380 2470 400
rect 2410 360 2430 380
rect 2450 360 2470 380
rect 2410 350 2470 360
rect 2520 325 2580 400
rect 2630 385 2690 400
rect 2520 305 2540 325
rect 2560 305 2580 325
rect 1970 270 2140 285
rect 1970 250 1990 270
rect 2010 250 2140 270
rect 1970 240 2140 250
rect 1970 230 2030 240
rect 2080 230 2140 240
rect 2190 270 2250 285
rect 2190 250 2210 270
rect 2230 250 2250 270
rect 2190 230 2250 250
rect 2300 270 2470 280
rect 2300 250 2375 270
rect 2395 250 2470 270
rect 2300 240 2470 250
rect 2300 230 2360 240
rect 2410 230 2470 240
rect 2520 230 2580 305
rect 2630 325 2690 335
rect 2630 305 2650 325
rect 2670 305 2690 325
rect 2630 230 2690 305
rect 2740 325 2800 400
rect 2740 305 2760 325
rect 2780 305 2800 325
rect 2740 230 2800 305
rect 2850 270 2910 400
rect 2850 250 2870 270
rect 2890 250 2910 270
rect 2850 230 2910 250
rect 0 65 60 80
rect 110 65 170 80
rect 220 65 280 80
rect 330 65 390 80
rect 440 65 500 80
rect 550 65 610 80
rect 660 65 720 80
rect 770 65 830 80
rect 880 65 940 80
rect 990 65 1050 80
rect 1100 65 1160 80
rect 1210 65 1270 80
rect 1320 65 1380 80
rect 1530 65 1590 80
rect 1640 65 1700 80
rect 1750 65 1810 80
rect 1860 65 1920 80
rect 1970 65 2030 80
rect 2080 65 2140 80
rect 2190 65 2250 80
rect 2300 65 2360 80
rect 2410 65 2470 80
rect 2520 65 2580 80
rect 2630 65 2690 80
rect 2740 65 2800 80
rect 2850 65 2910 80
<< polycont >>
rect 20 1455 40 1475
rect 130 1400 150 1420
rect 240 1400 260 1420
rect 515 1455 535 1475
rect 680 1455 700 1475
rect 900 1455 920 1475
rect 350 1400 370 1420
rect 460 1345 480 1365
rect 570 1345 590 1365
rect 1120 1400 1140 1420
rect 1770 1400 1790 1420
rect 1990 1455 2010 1475
rect 2210 1455 2230 1475
rect 2375 1455 2395 1475
rect 2540 1400 2560 1420
rect 2320 1345 2340 1365
rect 2430 1345 2450 1365
rect 2650 1400 2670 1420
rect 2760 1400 2780 1420
rect 2870 1455 2890 1475
rect 240 1125 260 1145
rect 680 1125 700 1145
rect 1010 1125 1030 1145
rect 1230 1125 1250 1145
rect 1340 1125 1360 1145
rect 1550 1125 1570 1145
rect 1660 1125 1680 1145
rect 1880 1125 1900 1145
rect 2210 1125 2230 1145
rect 2650 1125 2670 1145
rect 240 570 260 590
rect 680 570 700 590
rect 1010 570 1030 590
rect 1230 570 1250 590
rect 1340 570 1360 590
rect 1550 570 1570 590
rect 1660 570 1680 590
rect 1880 570 1900 590
rect 2210 570 2230 590
rect 2650 570 2670 590
rect 20 250 40 270
rect 130 305 150 325
rect 240 305 260 325
rect 460 360 480 380
rect 570 360 590 380
rect 350 305 370 325
rect 515 250 535 270
rect 680 250 700 270
rect 900 250 920 270
rect 1120 305 1140 325
rect 1230 250 1250 270
rect 1770 305 1790 325
rect 1660 250 1680 270
rect 2320 360 2340 380
rect 2430 360 2450 380
rect 2540 305 2560 325
rect 1990 250 2010 270
rect 2210 250 2230 270
rect 2375 250 2395 270
rect 2650 305 2670 325
rect 2760 305 2780 325
rect 2870 250 2890 270
<< locali >>
rect -215 1690 -175 1700
rect -215 1670 -205 1690
rect -185 1670 -175 1690
rect -215 535 -175 1670
rect 65 1690 105 1700
rect 65 1670 75 1690
rect 95 1670 105 1690
rect -95 1635 -5 1645
rect -95 1515 -85 1635
rect -65 1515 -35 1635
rect -15 1515 -5 1635
rect -95 1485 -5 1515
rect 65 1635 105 1670
rect 285 1690 325 1700
rect 285 1670 295 1690
rect 315 1670 325 1690
rect 65 1515 75 1635
rect 95 1515 105 1635
rect 65 1505 105 1515
rect 175 1635 215 1645
rect 175 1515 185 1635
rect 205 1515 215 1635
rect -95 1475 50 1485
rect -95 1455 20 1475
rect 40 1455 50 1475
rect -95 1445 50 1455
rect 175 1480 215 1515
rect 285 1635 325 1670
rect 2585 1690 2625 1700
rect 2585 1670 2595 1690
rect 2615 1670 2625 1690
rect 285 1515 295 1635
rect 315 1515 325 1635
rect 285 1505 325 1515
rect 395 1635 435 1645
rect 395 1515 405 1635
rect 425 1515 435 1635
rect 395 1505 435 1515
rect 505 1635 545 1645
rect 505 1515 515 1635
rect 535 1515 545 1635
rect 395 1480 430 1505
rect 175 1450 430 1480
rect -95 1305 -5 1445
rect 120 1420 270 1430
rect 120 1400 130 1420
rect 150 1400 185 1420
rect 205 1400 240 1420
rect 260 1400 270 1420
rect 120 1390 270 1400
rect 340 1420 380 1430
rect 340 1400 350 1420
rect 370 1400 380 1420
rect 340 1390 380 1400
rect -215 515 -205 535
rect -185 515 -175 535
rect -215 505 -175 515
rect -155 1205 -115 1215
rect -155 1185 -145 1205
rect -125 1185 -115 1205
rect -155 60 -115 1185
rect -95 1185 -85 1305
rect -65 1185 -35 1305
rect -15 1185 -5 1305
rect -95 1175 -5 1185
rect 65 1305 105 1315
rect 65 1185 75 1305
rect 95 1185 105 1305
rect 65 1175 105 1185
rect 175 1305 215 1390
rect 400 1315 430 1450
rect 505 1475 545 1515
rect 615 1635 655 1645
rect 615 1515 625 1635
rect 645 1515 655 1635
rect 615 1505 655 1515
rect 725 1635 765 1645
rect 725 1515 735 1635
rect 755 1535 765 1635
rect 945 1635 985 1645
rect 755 1515 870 1535
rect 725 1505 870 1515
rect 945 1515 955 1635
rect 975 1515 985 1635
rect 945 1505 985 1515
rect 1055 1635 1095 1645
rect 1055 1515 1065 1635
rect 1085 1515 1095 1635
rect 1055 1505 1095 1515
rect 1165 1635 1205 1645
rect 1165 1515 1175 1635
rect 1195 1515 1205 1635
rect 1165 1505 1205 1515
rect 1275 1635 1315 1645
rect 1275 1515 1285 1635
rect 1305 1515 1315 1635
rect 1275 1505 1315 1515
rect 1385 1635 1525 1645
rect 1385 1515 1395 1635
rect 1415 1515 1445 1635
rect 1465 1515 1495 1635
rect 1515 1515 1525 1635
rect 505 1455 515 1475
rect 535 1455 545 1475
rect 505 1445 545 1455
rect 450 1420 490 1430
rect 450 1400 460 1420
rect 480 1400 490 1420
rect 450 1365 490 1400
rect 450 1345 460 1365
rect 480 1345 490 1365
rect 450 1335 490 1345
rect 510 1315 540 1445
rect 560 1420 600 1430
rect 560 1400 570 1420
rect 590 1400 600 1420
rect 560 1365 600 1400
rect 560 1345 570 1365
rect 590 1345 600 1365
rect 560 1335 600 1345
rect 620 1315 650 1505
rect 670 1480 710 1485
rect 670 1475 815 1480
rect 670 1455 680 1475
rect 700 1455 815 1475
rect 670 1450 815 1455
rect 670 1445 710 1450
rect 175 1185 185 1305
rect 205 1185 215 1305
rect 175 1175 215 1185
rect 285 1305 325 1315
rect 285 1185 295 1305
rect 315 1185 325 1305
rect 285 1175 325 1185
rect 395 1305 435 1315
rect 395 1185 405 1305
rect 425 1185 435 1305
rect 395 1175 435 1185
rect 505 1305 545 1315
rect 505 1185 515 1305
rect 535 1185 545 1305
rect 505 1175 545 1185
rect 615 1305 655 1315
rect 615 1185 625 1305
rect 645 1185 655 1305
rect 615 1175 655 1185
rect 725 1305 765 1315
rect 725 1185 735 1305
rect 755 1185 765 1305
rect 725 1175 765 1185
rect 70 875 100 1175
rect 180 1095 210 1175
rect 230 1145 270 1155
rect 230 1125 240 1145
rect 260 1125 270 1145
rect 230 1115 270 1125
rect 290 1095 320 1175
rect 670 1150 710 1155
rect 565 1145 710 1150
rect 565 1125 680 1145
rect 700 1125 710 1145
rect 565 1120 710 1125
rect 120 1085 160 1095
rect 120 1065 130 1085
rect 150 1065 160 1085
rect 180 1065 265 1095
rect 120 1055 160 1065
rect 125 1030 155 1055
rect 235 1030 265 1065
rect 285 1085 325 1095
rect 285 1065 295 1085
rect 315 1065 325 1085
rect 285 1055 325 1065
rect 125 1000 210 1030
rect 235 1000 320 1030
rect 65 865 105 875
rect 65 845 75 865
rect 95 845 105 865
rect 65 835 105 845
rect 65 645 105 655
rect 65 625 75 645
rect 95 625 105 645
rect -95 535 -5 545
rect -95 415 -85 535
rect -65 415 -35 535
rect -15 415 -5 535
rect -95 280 -5 415
rect 65 535 105 625
rect 180 545 210 1000
rect 230 590 270 600
rect 230 570 240 590
rect 260 570 270 590
rect 230 560 270 570
rect 290 545 320 1000
rect 565 765 595 1120
rect 670 1115 710 1120
rect 730 1095 760 1175
rect 620 1065 760 1095
rect 785 1090 815 1450
rect 840 1150 870 1505
rect 890 1475 930 1485
rect 890 1455 900 1475
rect 920 1455 930 1475
rect 890 1445 930 1455
rect 950 1370 980 1505
rect 895 1340 980 1370
rect 1060 1370 1090 1505
rect 1110 1420 1150 1430
rect 1110 1400 1120 1420
rect 1140 1400 1150 1420
rect 1110 1390 1150 1400
rect 1060 1340 1145 1370
rect 835 1140 875 1150
rect 835 1120 845 1140
rect 865 1120 875 1140
rect 835 1110 875 1120
rect 560 755 600 765
rect 560 735 570 755
rect 590 735 600 755
rect 560 725 600 735
rect 620 655 650 1065
rect 785 1060 870 1090
rect 725 1030 765 1040
rect 725 1010 735 1030
rect 755 1010 765 1030
rect 725 1000 765 1010
rect 670 975 710 985
rect 670 955 680 975
rect 700 955 710 975
rect 670 945 710 955
rect 615 645 655 655
rect 615 625 625 645
rect 645 625 655 645
rect 615 615 655 625
rect 675 600 705 945
rect 670 590 710 600
rect 670 570 680 590
rect 700 570 710 590
rect 670 560 710 570
rect 730 545 760 1000
rect 840 985 870 1060
rect 835 975 875 985
rect 835 955 845 975
rect 865 955 875 975
rect 835 945 875 955
rect 895 930 925 1340
rect 945 1305 985 1315
rect 945 1185 955 1305
rect 975 1185 985 1305
rect 945 1175 985 1185
rect 1055 1305 1095 1315
rect 1055 1185 1065 1305
rect 1085 1185 1095 1305
rect 1055 1175 1095 1185
rect 950 1150 980 1175
rect 1000 1150 1040 1155
rect 950 1145 1040 1150
rect 950 1125 1010 1145
rect 1030 1125 1040 1145
rect 950 1120 1040 1125
rect 890 920 930 930
rect 890 900 900 920
rect 920 900 930 920
rect 890 890 930 900
rect 835 865 875 875
rect 835 845 845 865
rect 865 845 875 865
rect 835 835 875 845
rect 780 755 820 765
rect 780 735 790 755
rect 810 735 820 755
rect 780 725 820 735
rect 65 415 75 535
rect 95 415 105 535
rect 65 405 105 415
rect 175 535 215 545
rect 175 415 185 535
rect 205 415 215 535
rect 175 335 215 415
rect 285 535 325 545
rect 285 415 295 535
rect 315 415 325 535
rect 285 405 325 415
rect 395 535 435 545
rect 395 415 405 535
rect 425 415 435 535
rect 395 405 435 415
rect 505 535 545 545
rect 505 415 515 535
rect 535 415 545 535
rect 505 405 545 415
rect 615 535 655 545
rect 615 415 625 535
rect 645 415 655 535
rect 615 405 655 415
rect 725 535 765 545
rect 725 415 735 535
rect 755 415 765 535
rect 725 405 765 415
rect 120 325 270 335
rect 120 305 130 325
rect 150 305 185 325
rect 205 305 240 325
rect 260 305 270 325
rect 120 295 270 305
rect 340 325 380 335
rect 340 305 350 325
rect 370 305 380 325
rect 340 295 380 305
rect -95 270 50 280
rect 400 275 430 405
rect 450 380 490 390
rect 450 360 460 380
rect 480 360 490 380
rect 450 325 490 360
rect 450 305 460 325
rect 480 305 490 325
rect 450 295 490 305
rect 510 280 540 405
rect 560 380 600 390
rect 560 360 570 380
rect 590 360 600 380
rect 560 325 600 360
rect 560 305 570 325
rect 590 305 600 325
rect 560 295 600 305
rect -95 250 20 270
rect 40 250 50 270
rect -95 240 50 250
rect 175 245 430 275
rect -95 215 -5 240
rect -95 95 -85 215
rect -65 95 -35 215
rect -15 95 -5 215
rect -95 85 -5 95
rect 65 215 105 225
rect 65 95 75 215
rect 95 95 105 215
rect -155 40 -145 60
rect -125 40 -115 60
rect -155 30 -115 40
rect 65 60 105 95
rect 175 215 215 245
rect 395 225 430 245
rect 505 270 545 280
rect 505 250 515 270
rect 535 250 545 270
rect 175 95 185 215
rect 205 95 215 215
rect 175 85 215 95
rect 285 215 325 225
rect 285 95 295 215
rect 315 95 325 215
rect 65 40 75 60
rect 95 40 105 60
rect 65 30 105 40
rect 285 60 325 95
rect 395 215 435 225
rect 395 95 405 215
rect 425 95 435 215
rect 395 85 435 95
rect 505 215 545 250
rect 620 225 650 405
rect 670 275 710 280
rect 785 275 815 725
rect 670 270 815 275
rect 670 250 680 270
rect 700 250 815 270
rect 670 245 815 250
rect 670 240 710 245
rect 840 225 870 835
rect 895 385 925 890
rect 950 595 980 1120
rect 1000 1115 1040 1120
rect 1000 1085 1040 1095
rect 1000 1065 1010 1085
rect 1030 1065 1040 1085
rect 1000 1055 1040 1065
rect 1005 710 1035 1055
rect 1060 875 1090 1175
rect 1115 1040 1145 1340
rect 1170 1315 1200 1505
rect 1280 1315 1310 1505
rect 1165 1305 1205 1315
rect 1165 1185 1175 1305
rect 1195 1185 1205 1305
rect 1165 1175 1205 1185
rect 1275 1305 1315 1315
rect 1275 1185 1285 1305
rect 1305 1185 1315 1305
rect 1275 1175 1315 1185
rect 1385 1305 1525 1515
rect 1595 1635 1635 1645
rect 1595 1515 1605 1635
rect 1625 1515 1635 1635
rect 1595 1505 1635 1515
rect 1705 1635 1745 1645
rect 1705 1515 1715 1635
rect 1735 1515 1745 1635
rect 1705 1505 1745 1515
rect 1815 1635 1855 1645
rect 1815 1515 1825 1635
rect 1845 1515 1855 1635
rect 1815 1505 1855 1515
rect 1925 1635 1965 1645
rect 1925 1515 1935 1635
rect 1955 1515 1965 1635
rect 2145 1635 2185 1645
rect 2145 1535 2155 1635
rect 1925 1505 1965 1515
rect 2040 1515 2155 1535
rect 2175 1515 2185 1635
rect 2040 1505 2185 1515
rect 2255 1635 2295 1645
rect 2255 1515 2265 1635
rect 2285 1515 2295 1635
rect 2255 1505 2295 1515
rect 2365 1635 2405 1645
rect 2365 1515 2375 1635
rect 2395 1515 2405 1635
rect 1600 1315 1630 1505
rect 1710 1315 1740 1505
rect 1760 1420 1800 1430
rect 1760 1400 1770 1420
rect 1790 1400 1800 1420
rect 1760 1390 1800 1400
rect 1820 1370 1850 1505
rect 1765 1340 1850 1370
rect 1930 1370 1960 1505
rect 1980 1475 2020 1485
rect 1980 1455 1990 1475
rect 2010 1455 2020 1475
rect 1980 1445 2020 1455
rect 1930 1340 2015 1370
rect 1385 1185 1395 1305
rect 1415 1185 1445 1305
rect 1465 1185 1495 1305
rect 1515 1185 1525 1305
rect 1385 1175 1525 1185
rect 1595 1305 1635 1315
rect 1595 1185 1605 1305
rect 1625 1185 1635 1305
rect 1595 1175 1635 1185
rect 1705 1305 1745 1315
rect 1705 1185 1715 1305
rect 1735 1185 1745 1305
rect 1705 1175 1745 1185
rect 1220 1145 1260 1155
rect 1220 1125 1230 1145
rect 1250 1125 1260 1145
rect 1220 1115 1260 1125
rect 1110 1030 1150 1040
rect 1110 1010 1120 1030
rect 1140 1010 1150 1030
rect 1110 1000 1150 1010
rect 1225 930 1255 1115
rect 1220 920 1260 930
rect 1220 900 1230 920
rect 1250 900 1260 920
rect 1220 890 1260 900
rect 1055 865 1095 875
rect 1055 845 1065 865
rect 1085 845 1095 865
rect 1055 835 1095 845
rect 1280 820 1310 1175
rect 1330 1145 1370 1155
rect 1330 1125 1340 1145
rect 1360 1125 1370 1145
rect 1330 1115 1370 1125
rect 1540 1145 1580 1155
rect 1540 1125 1550 1145
rect 1570 1125 1580 1145
rect 1540 1115 1580 1125
rect 1335 930 1365 1115
rect 1545 930 1575 1115
rect 1330 920 1370 930
rect 1330 900 1340 920
rect 1360 900 1370 920
rect 1330 890 1370 900
rect 1540 920 1580 930
rect 1540 900 1550 920
rect 1570 900 1580 920
rect 1540 890 1580 900
rect 1275 810 1315 820
rect 1275 790 1285 810
rect 1305 790 1315 810
rect 1275 780 1315 790
rect 1000 700 1040 710
rect 1000 680 1010 700
rect 1030 680 1040 700
rect 1000 670 1040 680
rect 1110 700 1150 710
rect 1110 680 1120 700
rect 1140 680 1150 700
rect 1110 670 1150 680
rect 1055 645 1095 655
rect 1055 625 1065 645
rect 1085 625 1095 645
rect 1055 615 1095 625
rect 1000 595 1040 600
rect 950 590 1040 595
rect 950 570 1010 590
rect 1030 570 1040 590
rect 950 565 1040 570
rect 950 545 980 565
rect 1000 560 1040 565
rect 1060 545 1090 615
rect 945 535 985 545
rect 945 415 955 535
rect 975 415 985 535
rect 945 405 985 415
rect 1055 535 1095 545
rect 1055 415 1065 535
rect 1085 415 1095 535
rect 1055 405 1095 415
rect 1115 385 1145 670
rect 1165 590 1260 600
rect 1165 570 1230 590
rect 1250 570 1260 590
rect 1165 560 1260 570
rect 1165 535 1205 560
rect 1280 545 1310 780
rect 1335 600 1365 890
rect 1545 600 1575 890
rect 1600 820 1630 1175
rect 1650 1145 1690 1155
rect 1650 1125 1660 1145
rect 1680 1125 1690 1145
rect 1650 1115 1690 1125
rect 1655 930 1685 1115
rect 1765 1040 1795 1340
rect 1815 1305 1855 1315
rect 1815 1185 1825 1305
rect 1845 1185 1855 1305
rect 1815 1175 1855 1185
rect 1925 1305 1965 1315
rect 1925 1185 1935 1305
rect 1955 1185 1965 1305
rect 1925 1175 1965 1185
rect 1760 1030 1800 1040
rect 1760 1010 1770 1030
rect 1790 1010 1800 1030
rect 1760 1000 1800 1010
rect 1650 920 1690 930
rect 1650 900 1660 920
rect 1680 900 1690 920
rect 1650 890 1690 900
rect 1820 875 1850 1175
rect 1870 1150 1910 1155
rect 1930 1150 1960 1175
rect 1870 1145 1960 1150
rect 1870 1125 1880 1145
rect 1900 1125 1960 1145
rect 1870 1120 1960 1125
rect 1870 1115 1910 1120
rect 1870 1085 1910 1095
rect 1870 1065 1880 1085
rect 1900 1065 1910 1085
rect 1870 1055 1910 1065
rect 1815 865 1855 875
rect 1815 845 1825 865
rect 1845 845 1855 865
rect 1815 835 1855 845
rect 1595 810 1635 820
rect 1595 790 1605 810
rect 1625 790 1635 810
rect 1595 780 1635 790
rect 1330 590 1370 600
rect 1330 570 1340 590
rect 1360 570 1370 590
rect 1330 560 1370 570
rect 1540 590 1580 600
rect 1540 570 1550 590
rect 1570 570 1580 590
rect 1540 560 1580 570
rect 1600 545 1630 780
rect 1875 710 1905 1055
rect 1760 700 1800 710
rect 1760 680 1770 700
rect 1790 680 1800 700
rect 1760 670 1800 680
rect 1870 700 1910 710
rect 1870 680 1880 700
rect 1900 680 1910 700
rect 1870 670 1910 680
rect 1650 590 1745 600
rect 1650 570 1660 590
rect 1680 570 1745 590
rect 1650 560 1745 570
rect 1165 415 1175 535
rect 1195 415 1205 535
rect 1165 405 1205 415
rect 1275 535 1315 545
rect 1275 415 1285 535
rect 1305 415 1315 535
rect 1275 405 1315 415
rect 1385 535 1525 545
rect 1385 415 1395 535
rect 1415 415 1445 535
rect 1465 415 1495 535
rect 1515 415 1525 535
rect 895 355 980 385
rect 890 270 930 280
rect 890 250 900 270
rect 920 250 930 270
rect 890 240 930 250
rect 950 225 980 355
rect 1060 355 1145 385
rect 1060 225 1090 355
rect 1110 325 1150 335
rect 1110 305 1120 325
rect 1140 305 1150 325
rect 1110 295 1150 305
rect 1170 280 1200 405
rect 1165 270 1260 280
rect 1165 250 1230 270
rect 1250 250 1260 270
rect 1165 240 1260 250
rect 505 95 515 215
rect 535 95 545 215
rect 505 85 545 95
rect 615 215 655 225
rect 615 95 625 215
rect 645 95 655 215
rect 615 85 655 95
rect 725 215 870 225
rect 725 95 735 215
rect 755 195 870 215
rect 945 215 985 225
rect 755 95 765 195
rect 725 85 765 95
rect 945 95 955 215
rect 975 95 985 215
rect 945 85 985 95
rect 1055 215 1095 225
rect 1055 95 1065 215
rect 1085 95 1095 215
rect 1055 85 1095 95
rect 1165 215 1205 240
rect 1280 225 1310 405
rect 1165 95 1175 215
rect 1195 95 1205 215
rect 1165 85 1205 95
rect 1275 215 1315 225
rect 1275 95 1285 215
rect 1305 95 1315 215
rect 1275 85 1315 95
rect 1385 215 1525 415
rect 1595 535 1635 545
rect 1595 415 1605 535
rect 1625 415 1635 535
rect 1595 405 1635 415
rect 1705 535 1745 560
rect 1705 415 1715 535
rect 1735 415 1745 535
rect 1705 405 1745 415
rect 1600 225 1630 405
rect 1710 280 1740 405
rect 1765 385 1795 670
rect 1815 645 1855 655
rect 1815 625 1825 645
rect 1845 625 1855 645
rect 1815 615 1855 625
rect 1820 545 1850 615
rect 1870 595 1910 600
rect 1930 595 1960 1120
rect 1985 930 2015 1340
rect 2040 1150 2070 1505
rect 2200 1480 2240 1485
rect 2095 1475 2240 1480
rect 2095 1455 2210 1475
rect 2230 1455 2240 1475
rect 2095 1450 2240 1455
rect 2035 1140 2075 1150
rect 2035 1120 2045 1140
rect 2065 1120 2075 1140
rect 2035 1110 2075 1120
rect 2095 1090 2125 1450
rect 2200 1445 2240 1450
rect 2260 1315 2290 1505
rect 2365 1475 2405 1515
rect 2475 1635 2515 1645
rect 2475 1515 2485 1635
rect 2505 1515 2515 1635
rect 2475 1505 2515 1515
rect 2585 1635 2625 1670
rect 2805 1690 2845 1700
rect 2805 1670 2815 1690
rect 2835 1670 2845 1690
rect 2585 1515 2595 1635
rect 2615 1515 2625 1635
rect 2585 1505 2625 1515
rect 2695 1635 2735 1645
rect 2695 1515 2705 1635
rect 2725 1515 2735 1635
rect 2365 1455 2375 1475
rect 2395 1455 2405 1475
rect 2365 1445 2405 1455
rect 2480 1480 2515 1505
rect 2695 1480 2735 1515
rect 2805 1635 2845 1670
rect 3085 1690 3125 1700
rect 3085 1670 3095 1690
rect 3115 1670 3125 1690
rect 2805 1515 2815 1635
rect 2835 1515 2845 1635
rect 2805 1505 2845 1515
rect 2915 1635 3005 1645
rect 2915 1515 2925 1635
rect 2945 1515 2975 1635
rect 2995 1515 3005 1635
rect 2915 1485 3005 1515
rect 2480 1450 2735 1480
rect 2860 1475 3005 1485
rect 2860 1455 2870 1475
rect 2890 1455 3005 1475
rect 2310 1420 2350 1430
rect 2310 1400 2320 1420
rect 2340 1400 2350 1420
rect 2310 1365 2350 1400
rect 2310 1345 2320 1365
rect 2340 1345 2350 1365
rect 2310 1335 2350 1345
rect 2370 1315 2400 1445
rect 2420 1420 2460 1430
rect 2420 1400 2430 1420
rect 2450 1400 2460 1420
rect 2420 1365 2460 1400
rect 2420 1345 2430 1365
rect 2450 1345 2460 1365
rect 2420 1335 2460 1345
rect 2480 1315 2510 1450
rect 2860 1445 3005 1455
rect 2530 1420 2570 1430
rect 2530 1400 2540 1420
rect 2560 1400 2570 1420
rect 2530 1390 2570 1400
rect 2640 1420 2790 1430
rect 2640 1400 2650 1420
rect 2670 1400 2705 1420
rect 2725 1400 2760 1420
rect 2780 1400 2790 1420
rect 2640 1390 2790 1400
rect 2145 1305 2185 1315
rect 2145 1185 2155 1305
rect 2175 1185 2185 1305
rect 2145 1175 2185 1185
rect 2255 1305 2295 1315
rect 2255 1185 2265 1305
rect 2285 1185 2295 1305
rect 2255 1175 2295 1185
rect 2365 1305 2405 1315
rect 2365 1185 2375 1305
rect 2395 1185 2405 1305
rect 2365 1175 2405 1185
rect 2475 1305 2515 1315
rect 2475 1185 2485 1305
rect 2505 1185 2515 1305
rect 2475 1175 2515 1185
rect 2585 1305 2625 1315
rect 2585 1185 2595 1305
rect 2615 1185 2625 1305
rect 2585 1175 2625 1185
rect 2695 1305 2735 1390
rect 2695 1185 2705 1305
rect 2725 1185 2735 1305
rect 2695 1175 2735 1185
rect 2805 1305 2845 1315
rect 2805 1185 2815 1305
rect 2835 1185 2845 1305
rect 2805 1175 2845 1185
rect 2915 1305 3005 1445
rect 2915 1185 2925 1305
rect 2945 1185 2975 1305
rect 2995 1185 3005 1305
rect 2915 1175 3005 1185
rect 3025 1205 3065 1215
rect 3025 1185 3035 1205
rect 3055 1185 3065 1205
rect 2040 1060 2125 1090
rect 2150 1095 2180 1175
rect 2200 1150 2240 1155
rect 2200 1145 2345 1150
rect 2200 1125 2210 1145
rect 2230 1125 2345 1145
rect 2200 1120 2345 1125
rect 2200 1115 2240 1120
rect 2150 1065 2290 1095
rect 2040 985 2070 1060
rect 2145 1030 2185 1040
rect 2145 1010 2155 1030
rect 2175 1010 2185 1030
rect 2145 1000 2185 1010
rect 2035 975 2075 985
rect 2035 955 2045 975
rect 2065 955 2075 975
rect 2035 945 2075 955
rect 1980 920 2020 930
rect 1980 900 1990 920
rect 2010 900 2020 920
rect 1980 890 2020 900
rect 1870 590 1960 595
rect 1870 570 1880 590
rect 1900 570 1960 590
rect 1870 565 1960 570
rect 1870 560 1910 565
rect 1930 545 1960 565
rect 1815 535 1855 545
rect 1815 415 1825 535
rect 1845 415 1855 535
rect 1815 405 1855 415
rect 1925 535 1965 545
rect 1925 415 1935 535
rect 1955 415 1965 535
rect 1925 405 1965 415
rect 1985 385 2015 890
rect 2035 865 2075 875
rect 2035 845 2045 865
rect 2065 845 2075 865
rect 2035 835 2075 845
rect 1765 355 1850 385
rect 1760 325 1800 335
rect 1760 305 1770 325
rect 1790 305 1800 325
rect 1760 295 1800 305
rect 1650 270 1745 280
rect 1650 250 1660 270
rect 1680 250 1745 270
rect 1650 240 1745 250
rect 1385 95 1395 215
rect 1415 95 1445 215
rect 1465 95 1495 215
rect 1515 95 1525 215
rect 1385 85 1525 95
rect 1595 215 1635 225
rect 1595 95 1605 215
rect 1625 95 1635 215
rect 1595 85 1635 95
rect 1705 215 1745 240
rect 1820 225 1850 355
rect 1930 355 2015 385
rect 1930 225 1960 355
rect 1980 270 2020 280
rect 1980 250 1990 270
rect 2010 250 2020 270
rect 1980 240 2020 250
rect 2040 225 2070 835
rect 2090 755 2130 765
rect 2090 735 2100 755
rect 2120 735 2130 755
rect 2090 725 2130 735
rect 2095 275 2125 725
rect 2150 545 2180 1000
rect 2200 975 2240 985
rect 2200 955 2210 975
rect 2230 955 2240 975
rect 2200 945 2240 955
rect 2205 600 2235 945
rect 2260 655 2290 1065
rect 2315 765 2345 1120
rect 2590 1095 2620 1175
rect 2640 1145 2680 1155
rect 2640 1125 2650 1145
rect 2670 1125 2680 1145
rect 2640 1115 2680 1125
rect 2700 1095 2730 1175
rect 2585 1085 2625 1095
rect 2585 1065 2595 1085
rect 2615 1065 2625 1085
rect 2585 1055 2625 1065
rect 2645 1065 2730 1095
rect 2750 1085 2790 1095
rect 2750 1065 2760 1085
rect 2780 1065 2790 1085
rect 2645 1030 2675 1065
rect 2750 1055 2790 1065
rect 2755 1030 2785 1055
rect 2590 1000 2675 1030
rect 2700 1000 2785 1030
rect 2310 755 2350 765
rect 2310 735 2320 755
rect 2340 735 2350 755
rect 2310 725 2350 735
rect 2255 645 2295 655
rect 2255 625 2265 645
rect 2285 625 2295 645
rect 2255 615 2295 625
rect 2200 590 2240 600
rect 2200 570 2210 590
rect 2230 570 2240 590
rect 2200 560 2240 570
rect 2590 545 2620 1000
rect 2640 590 2680 600
rect 2640 570 2650 590
rect 2670 570 2680 590
rect 2640 560 2680 570
rect 2700 545 2730 1000
rect 2810 875 2840 1175
rect 2805 865 2845 875
rect 2805 845 2815 865
rect 2835 845 2845 865
rect 2805 835 2845 845
rect 2805 645 2845 655
rect 2805 625 2815 645
rect 2835 625 2845 645
rect 2145 535 2185 545
rect 2145 415 2155 535
rect 2175 415 2185 535
rect 2145 405 2185 415
rect 2255 535 2295 545
rect 2255 415 2265 535
rect 2285 415 2295 535
rect 2255 405 2295 415
rect 2365 535 2405 545
rect 2365 415 2375 535
rect 2395 415 2405 535
rect 2365 405 2405 415
rect 2475 535 2515 545
rect 2475 415 2485 535
rect 2505 415 2515 535
rect 2475 405 2515 415
rect 2585 535 2625 545
rect 2585 415 2595 535
rect 2615 415 2625 535
rect 2585 405 2625 415
rect 2695 535 2735 545
rect 2695 415 2705 535
rect 2725 415 2735 535
rect 2200 275 2240 280
rect 2095 270 2240 275
rect 2095 250 2210 270
rect 2230 250 2240 270
rect 2095 245 2240 250
rect 2200 240 2240 245
rect 2260 225 2290 405
rect 2310 380 2350 390
rect 2310 360 2320 380
rect 2340 360 2350 380
rect 2310 325 2350 360
rect 2310 305 2320 325
rect 2340 305 2350 325
rect 2310 295 2350 305
rect 2370 280 2400 405
rect 2420 380 2460 390
rect 2420 360 2430 380
rect 2450 360 2460 380
rect 2420 325 2460 360
rect 2420 305 2430 325
rect 2450 305 2460 325
rect 2420 295 2460 305
rect 2365 270 2405 280
rect 2365 250 2375 270
rect 2395 250 2405 270
rect 1705 95 1715 215
rect 1735 95 1745 215
rect 1705 85 1745 95
rect 1815 215 1855 225
rect 1815 95 1825 215
rect 1845 95 1855 215
rect 1815 85 1855 95
rect 1925 215 1965 225
rect 1925 95 1935 215
rect 1955 95 1965 215
rect 2040 215 2185 225
rect 2040 195 2155 215
rect 1925 85 1965 95
rect 2145 95 2155 195
rect 2175 95 2185 215
rect 2145 85 2185 95
rect 2255 215 2295 225
rect 2255 95 2265 215
rect 2285 95 2295 215
rect 2255 85 2295 95
rect 2365 215 2405 250
rect 2480 275 2510 405
rect 2695 335 2735 415
rect 2805 535 2845 625
rect 2805 415 2815 535
rect 2835 415 2845 535
rect 2805 405 2845 415
rect 2915 535 3005 545
rect 2915 415 2925 535
rect 2945 415 2975 535
rect 2995 415 3005 535
rect 2530 325 2570 335
rect 2530 305 2540 325
rect 2560 305 2570 325
rect 2530 295 2570 305
rect 2640 325 2790 335
rect 2640 305 2650 325
rect 2670 305 2705 325
rect 2725 305 2760 325
rect 2780 305 2790 325
rect 2640 295 2790 305
rect 2915 280 3005 415
rect 2480 245 2735 275
rect 2480 225 2515 245
rect 2365 95 2375 215
rect 2395 95 2405 215
rect 2365 85 2405 95
rect 2475 215 2515 225
rect 2475 95 2485 215
rect 2505 95 2515 215
rect 2475 85 2515 95
rect 2585 215 2625 225
rect 2585 95 2595 215
rect 2615 95 2625 215
rect 285 40 295 60
rect 315 40 325 60
rect 285 30 325 40
rect 2585 60 2625 95
rect 2695 215 2735 245
rect 2860 270 3005 280
rect 2860 250 2870 270
rect 2890 250 3005 270
rect 2860 240 3005 250
rect 2695 95 2705 215
rect 2725 95 2735 215
rect 2695 85 2735 95
rect 2805 215 2845 225
rect 2805 95 2815 215
rect 2835 95 2845 215
rect 2585 40 2595 60
rect 2615 40 2625 60
rect 2585 30 2625 40
rect 2805 60 2845 95
rect 2915 215 3005 240
rect 2915 95 2925 215
rect 2945 95 2975 215
rect 2995 95 3005 215
rect 2915 85 3005 95
rect 2805 40 2815 60
rect 2835 40 2845 60
rect 2805 30 2845 40
rect 3025 60 3065 1185
rect 3085 535 3125 1670
rect 3085 515 3095 535
rect 3115 515 3125 535
rect 3085 505 3125 515
rect 3145 975 3185 985
rect 3145 955 3155 975
rect 3175 955 3185 975
rect 3145 365 3185 955
rect 3145 345 3155 365
rect 3175 345 3185 365
rect 3145 335 3185 345
rect 3205 755 3245 765
rect 3205 735 3215 755
rect 3235 735 3245 755
rect 3205 305 3245 735
rect 3205 285 3215 305
rect 3235 285 3245 305
rect 3205 275 3245 285
rect 3025 40 3035 60
rect 3055 40 3065 60
rect 3025 30 3065 40
<< viali >>
rect -205 1670 -185 1690
rect 75 1670 95 1690
rect -85 1515 -65 1635
rect -35 1515 -15 1635
rect 295 1670 315 1690
rect 2595 1670 2615 1690
rect 515 1515 535 1635
rect 130 1400 150 1420
rect 185 1400 205 1420
rect 240 1400 260 1420
rect 350 1400 370 1420
rect -205 515 -185 535
rect -145 1185 -125 1205
rect -85 1185 -65 1305
rect -35 1185 -15 1305
rect 1175 1515 1195 1635
rect 1395 1515 1415 1635
rect 1445 1515 1465 1635
rect 1495 1515 1515 1635
rect 460 1400 480 1420
rect 570 1400 590 1420
rect 515 1185 535 1305
rect 240 1125 260 1145
rect 130 1065 150 1085
rect 295 1065 315 1085
rect 75 845 95 865
rect 75 625 95 645
rect -85 415 -65 535
rect -35 415 -15 535
rect 240 570 260 590
rect 900 1455 920 1475
rect 1120 1400 1140 1420
rect 845 1120 865 1140
rect 570 735 590 755
rect 735 1010 755 1030
rect 680 955 700 975
rect 625 625 645 645
rect 845 955 865 975
rect 900 900 920 920
rect 845 845 865 865
rect 790 735 810 755
rect 515 415 535 535
rect 130 305 150 325
rect 185 305 205 325
rect 240 305 260 325
rect 350 305 370 325
rect 460 305 480 325
rect 570 305 590 325
rect -85 95 -65 215
rect -35 95 -15 215
rect -145 40 -125 60
rect 75 40 95 60
rect 1010 1065 1030 1085
rect 1175 1185 1195 1305
rect 1715 1515 1735 1635
rect 2375 1515 2395 1635
rect 1770 1400 1790 1420
rect 1990 1455 2010 1475
rect 1395 1185 1415 1305
rect 1445 1185 1465 1305
rect 1495 1185 1515 1305
rect 1715 1185 1735 1305
rect 1120 1010 1140 1030
rect 1230 900 1250 920
rect 1065 845 1085 865
rect 1340 900 1360 920
rect 1550 900 1570 920
rect 1285 790 1305 810
rect 1010 680 1030 700
rect 1120 680 1140 700
rect 1065 625 1085 645
rect 1770 1010 1790 1030
rect 1660 900 1680 920
rect 1880 1065 1900 1085
rect 1825 845 1845 865
rect 1605 790 1625 810
rect 1770 680 1790 700
rect 1880 680 1900 700
rect 1175 415 1195 535
rect 1395 415 1415 535
rect 1445 415 1465 535
rect 1495 415 1515 535
rect 900 250 920 270
rect 1120 305 1140 325
rect 515 95 535 215
rect 1175 95 1195 215
rect 1715 415 1735 535
rect 1825 625 1845 645
rect 2045 1120 2065 1140
rect 2815 1670 2835 1690
rect 3095 1670 3115 1690
rect 2925 1515 2945 1635
rect 2975 1515 2995 1635
rect 2320 1400 2340 1420
rect 2430 1400 2450 1420
rect 2540 1400 2560 1420
rect 2650 1400 2670 1420
rect 2705 1400 2725 1420
rect 2760 1400 2780 1420
rect 2375 1185 2395 1305
rect 2925 1185 2945 1305
rect 2975 1185 2995 1305
rect 3035 1185 3055 1205
rect 2155 1010 2175 1030
rect 2045 955 2065 975
rect 1990 900 2010 920
rect 2045 845 2065 865
rect 1770 305 1790 325
rect 1395 95 1415 215
rect 1445 95 1465 215
rect 1495 95 1515 215
rect 1990 250 2010 270
rect 2100 735 2120 755
rect 2210 955 2230 975
rect 2650 1125 2670 1145
rect 2595 1065 2615 1085
rect 2760 1065 2780 1085
rect 2320 735 2340 755
rect 2265 625 2285 645
rect 2650 570 2670 590
rect 2815 845 2835 865
rect 2815 625 2835 645
rect 2375 415 2395 535
rect 2320 305 2340 325
rect 2430 305 2450 325
rect 1715 95 1735 215
rect 2925 415 2945 535
rect 2975 415 2995 535
rect 2540 305 2560 325
rect 2650 305 2670 325
rect 2705 305 2725 325
rect 2760 305 2780 325
rect 2375 95 2395 215
rect 295 40 315 60
rect 2595 40 2615 60
rect 2925 95 2945 215
rect 2975 95 2995 215
rect 2815 40 2835 60
rect 3095 515 3115 535
rect 3155 955 3175 975
rect 3155 345 3175 365
rect 3215 735 3235 755
rect 3215 285 3235 305
rect 3035 40 3055 60
<< metal1 >>
rect -215 1690 3125 1700
rect -215 1670 -205 1690
rect -185 1670 75 1690
rect 95 1670 295 1690
rect 315 1670 2595 1690
rect 2615 1670 2815 1690
rect 2835 1670 3095 1690
rect 3115 1670 3125 1690
rect -215 1660 3125 1670
rect -230 1635 3140 1645
rect -230 1515 -85 1635
rect -65 1515 -35 1635
rect -15 1515 515 1635
rect 535 1515 1175 1635
rect 1195 1515 1395 1635
rect 1415 1515 1445 1635
rect 1465 1515 1495 1635
rect 1515 1515 1715 1635
rect 1735 1515 2375 1635
rect 2395 1515 2925 1635
rect 2945 1515 2975 1635
rect 2995 1515 3140 1635
rect -230 1505 3140 1515
rect -230 1315 -5 1505
rect 890 1475 930 1505
rect 890 1455 900 1475
rect 920 1455 930 1475
rect 890 1445 930 1455
rect 1980 1475 2020 1505
rect 1980 1455 1990 1475
rect 2010 1455 2020 1475
rect 1980 1445 2020 1455
rect 120 1420 2790 1430
rect 120 1400 130 1420
rect 150 1400 185 1420
rect 205 1400 240 1420
rect 260 1400 350 1420
rect 370 1400 460 1420
rect 480 1400 570 1420
rect 590 1400 1120 1420
rect 1140 1400 1770 1420
rect 1790 1400 2320 1420
rect 2340 1400 2430 1420
rect 2450 1400 2540 1420
rect 2560 1400 2650 1420
rect 2670 1400 2705 1420
rect 2725 1400 2760 1420
rect 2780 1400 2790 1420
rect 120 1390 2790 1400
rect 2915 1315 3140 1505
rect -230 1305 3140 1315
rect -230 1205 -85 1305
rect -230 1185 -145 1205
rect -125 1185 -85 1205
rect -65 1185 -35 1305
rect -15 1185 515 1305
rect 535 1185 1175 1305
rect 1195 1185 1395 1305
rect 1415 1185 1445 1305
rect 1465 1185 1495 1305
rect 1515 1185 1715 1305
rect 1735 1185 2375 1305
rect 2395 1185 2925 1305
rect 2945 1185 2975 1305
rect 2995 1205 3140 1305
rect 2995 1185 3035 1205
rect 3055 1185 3140 1205
rect -230 1175 3140 1185
rect 230 1145 270 1175
rect 230 1125 240 1145
rect 260 1125 270 1145
rect 230 1115 270 1125
rect 835 1140 875 1150
rect 835 1120 845 1140
rect 865 1120 875 1140
rect 835 1095 875 1120
rect 2035 1140 2075 1150
rect 2035 1120 2045 1140
rect 2065 1120 2075 1140
rect 2035 1095 2075 1120
rect 2640 1145 2680 1175
rect 2640 1125 2650 1145
rect 2670 1125 2680 1145
rect 2640 1115 2680 1125
rect 3175 1100 3245 1105
rect 120 1085 325 1095
rect 120 1065 130 1085
rect 150 1065 295 1085
rect 315 1065 325 1085
rect 120 1055 325 1065
rect 835 1085 1040 1095
rect 835 1065 1010 1085
rect 1030 1065 1040 1085
rect 835 1055 1040 1065
rect 1870 1085 2075 1095
rect 1870 1065 1880 1085
rect 1900 1065 2075 1085
rect 1870 1055 2075 1065
rect 2585 1085 2790 1095
rect 2585 1065 2595 1085
rect 2615 1065 2760 1085
rect 2780 1065 2790 1085
rect 2585 1055 2790 1065
rect 3175 1060 3180 1100
rect 3220 1060 3245 1100
rect 3175 1055 3245 1060
rect -100 1030 3010 1040
rect -100 1010 735 1030
rect 755 1010 1120 1030
rect 1140 1010 1770 1030
rect 1790 1010 2155 1030
rect 2175 1010 3010 1030
rect -100 1000 3010 1010
rect -230 975 3185 985
rect -230 955 680 975
rect 700 955 845 975
rect 865 955 2045 975
rect 2065 955 2210 975
rect 2230 955 3155 975
rect 3175 955 3185 975
rect -230 945 3185 955
rect 3205 930 3245 1055
rect -100 920 3245 930
rect -100 900 900 920
rect 920 900 1230 920
rect 1250 900 1340 920
rect 1360 900 1550 920
rect 1570 900 1660 920
rect 1680 900 1990 920
rect 2010 900 3245 920
rect -100 890 3245 900
rect -100 865 3015 875
rect -100 845 75 865
rect 95 845 845 865
rect 865 845 1065 865
rect 1085 845 1825 865
rect 1845 845 2045 865
rect 2065 845 2815 865
rect 2835 845 3015 865
rect -100 835 3015 845
rect 3205 870 3255 875
rect 3205 830 3210 870
rect 3250 830 3255 870
rect 3205 820 3255 830
rect -230 810 3255 820
rect -230 790 1285 810
rect 1305 790 1605 810
rect 1625 790 3255 810
rect -230 780 3255 790
rect -230 755 3245 765
rect -230 735 570 755
rect 590 735 790 755
rect 810 735 2100 755
rect 2120 735 2320 755
rect 2340 735 3215 755
rect 3235 735 3245 755
rect -230 725 3245 735
rect -100 700 3010 710
rect -100 680 1010 700
rect 1030 680 1120 700
rect 1140 680 1770 700
rect 1790 680 1880 700
rect 1900 680 3010 700
rect -100 670 3010 680
rect -100 645 3010 655
rect -100 625 75 645
rect 95 625 625 645
rect 645 625 1065 645
rect 1085 625 1825 645
rect 1845 625 2265 645
rect 2285 625 2815 645
rect 2835 625 3010 645
rect -100 615 3010 625
rect 230 590 270 600
rect 230 570 240 590
rect 260 570 270 590
rect -230 545 -5 560
rect 230 545 270 570
rect 2640 590 2680 600
rect 2640 570 2650 590
rect 2670 570 2680 590
rect 2640 545 2680 570
rect 2915 545 3125 560
rect -230 535 3125 545
rect -230 515 -205 535
rect -185 515 -85 535
rect -230 415 -85 515
rect -65 415 -35 535
rect -15 415 515 535
rect 535 415 1175 535
rect 1195 415 1395 535
rect 1415 415 1445 535
rect 1465 415 1495 535
rect 1515 415 1715 535
rect 1735 415 2375 535
rect 2395 415 2925 535
rect 2945 415 2975 535
rect 2995 515 3095 535
rect 3115 515 3125 535
rect 2995 415 3125 515
rect 5340 470 5390 475
rect 5340 430 5345 470
rect 5385 465 5390 470
rect 5385 430 5425 465
rect 5340 425 5425 430
rect -230 405 3125 415
rect -230 225 -5 405
rect 120 325 2790 335
rect 120 305 130 325
rect 150 305 185 325
rect 205 305 240 325
rect 260 305 350 325
rect 370 305 460 325
rect 480 305 570 325
rect 590 305 1120 325
rect 1140 305 1770 325
rect 1790 305 2320 325
rect 2340 305 2430 325
rect 2450 305 2540 325
rect 2560 305 2650 325
rect 2670 305 2705 325
rect 2725 305 2760 325
rect 2780 305 2790 325
rect 120 295 2790 305
rect 890 270 930 280
rect 890 250 900 270
rect 920 250 930 270
rect 890 225 930 250
rect 1980 270 2020 280
rect 1980 250 1990 270
rect 2010 250 2020 270
rect 1980 225 2020 250
rect 2915 225 3125 405
rect 3145 365 5425 375
rect 3145 345 3155 365
rect 3175 345 5425 365
rect 3145 335 5425 345
rect 3165 305 5425 315
rect 3165 285 3215 305
rect 3235 285 5425 305
rect 3165 275 5425 285
rect -230 215 3125 225
rect -230 95 -85 215
rect -65 95 -35 215
rect -15 95 515 215
rect 535 95 1175 215
rect 1195 95 1395 215
rect 1415 95 1445 215
rect 1465 95 1495 215
rect 1515 95 1715 215
rect 1735 95 2375 215
rect 2395 95 2925 215
rect 2945 95 2975 215
rect 2995 95 3125 215
rect -230 85 3125 95
rect -155 60 3065 70
rect -155 40 -145 60
rect -125 40 75 60
rect 95 40 295 60
rect 315 40 2595 60
rect 2615 40 2815 60
rect 2835 40 3035 60
rect 3055 40 3065 60
rect -155 30 3065 40
<< via1 >>
rect 3180 1060 3220 1100
rect 3210 830 3250 870
rect 5345 430 5385 470
<< metal2 >>
rect 3175 1100 3225 1105
rect 3175 1060 3180 1100
rect 3220 1060 3225 1100
rect 3175 1055 3225 1060
rect 3205 870 3255 875
rect 3205 830 3210 870
rect 3250 830 3255 870
rect 3205 825 3255 830
rect 5340 470 5390 475
rect 5340 430 5345 470
rect 5385 430 5390 470
rect 5340 425 5390 430
<< via2 >>
rect 3180 1060 3220 1100
rect 3210 830 3250 870
rect 5345 430 5385 470
<< metal3 >>
rect 3175 1100 3225 1105
rect 3175 1060 3180 1100
rect 3220 1060 3225 1100
rect 3175 1055 3225 1060
rect 3265 875 5295 1655
rect 3205 870 5295 875
rect 3205 830 3210 870
rect 3250 830 5295 870
rect 3205 825 5295 830
rect 3265 475 5295 825
rect 3265 470 5390 475
rect 3265 430 5345 470
rect 5385 430 5390 470
rect 3265 425 5390 430
<< via3 >>
rect 3180 1060 3220 1100
<< mimcap >>
rect 3280 1095 5280 1640
rect 3280 1060 3290 1095
rect 3325 1060 5280 1095
rect 3280 440 5280 1060
<< mimcapcontact >>
rect 3290 1060 3325 1095
<< metal4 >>
rect 3175 1100 3225 1105
rect 3175 1060 3180 1100
rect 3220 1095 3330 1100
rect 3220 1060 3290 1095
rect 3325 1060 3330 1095
rect 3175 1055 3330 1060
<< labels >>
rlabel metal1 -230 1175 -215 1645 7 vdd
port 4 w
rlabel metal1 -230 85 -215 560 7 gnd
port 5 w
rlabel ndiff 830 80 880 230 5 net16
rlabel ndiff 830 400 880 550 5 net15
rlabel pdiff 830 1170 880 1320 1 net14
rlabel pdiff 830 1500 880 1650 1 net13
rlabel pdiff 2030 1500 2080 1650 1 net22
rlabel locali 1055 1505 1095 1645 1 net3
rlabel locali 1055 1175 1095 1315 1 net4
rlabel locali 1055 405 1095 545 5 net7
rlabel locali 1055 85 1095 225 5 net6
rlabel locali 945 1175 985 1315 1 net5
rlabel locali 945 1505 985 1645 1 net2
rlabel metal1 120 1390 160 1430 7 net10
rlabel metal1 120 295 160 335 7 net9
rlabel locali 175 1505 215 1645 1 net12
rlabel locali 175 85 215 225 5 net1
rlabel locali 615 1505 655 1645 5 net11
rlabel locali 615 405 655 545 1 net8
rlabel metal1 -230 945 -215 985 7 v1
port 1 w
rlabel metal1 -230 725 -215 765 7 v2
port 2 w
rlabel metal1 -230 780 -215 820 7 vout
port 3 w
<< end >>
