* SPICE3 file created from error_amp.ext - technology: sky130A

.subckt k_res VSUBS a_n10_780# a_1270_n10#
X0 a_n10_n10# a_310_780# VSUBS sky130_fd_pr__res_xhigh_po w=0.35 l=1.75
X1 a_n10_n10# a_n10_780# VSUBS sky130_fd_pr__res_xhigh_po w=0.35 l=1.75
X2 a_630_n10# a_310_780# VSUBS sky130_fd_pr__res_xhigh_po w=0.35 l=1.75
X3 a_1270_n10# a_950_780# VSUBS sky130_fd_pr__res_xhigh_po w=0.35 l=1.75
X4 a_630_n10# a_950_780# VSUBS sky130_fd_pr__res_xhigh_po w=0.35 l=1.75
.ends

.subckt opamp v1 v2 vout vdd gnd
X0 vout net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=3e+12p pd=1.6e+07u as=1.2e+13p ps=6.4e+07u w=1.5e+06u l=600000u
X1 net7 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=3e+12p pd=1.6e+07u as=0p ps=0u w=1.5e+06u l=600000u
X2 net2 a_3720_130# net3 vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X3 net6 net5 net2 gnd sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X4 gnd net9 net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X5 gnd net2 vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X6 net7 vdd a_4060_2340# vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X7 vdd net10 net12 vdd sky130_fd_pr__pfet_01v8 ad=1.2e+13p pd=6.4e+07u as=2.25e+12p ps=1.2e+07u w=1.5e+06u l=600000u
X8 vdd vdd net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.6e+07u w=1.5e+06u l=600000u
X9 a_4060_160# gnd net2 gnd sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X10 net3 gnd a_4060_800# gnd sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X11 gnd net9 a_4500_160# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X12 net10 gnd net9 gnd sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X13 net4 net10 net10 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X14 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.6e+07u as=0p ps=0u w=1.5e+06u l=600000u
X15 net5 vdd net14 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X16 vdd net10 a_4500_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X17 gnd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=7.5e+12p pd=4e+07u as=0p ps=0u w=1.5e+06u l=600000u
X18 gnd gnd net1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=2.25e+12p ps=1.2e+07u w=1.5e+06u l=600000u
X19 net7 gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X20 net9 gnd net10 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X21 gnd gnd net7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X22 net22 vdd net2 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X23 net12 net10 gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X24 net3 v1 net8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X25 vdd net10 net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X26 a_4500_2340# v2 net7 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X27 net4 net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X28 net2 gnd net16 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X29 vout gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X30 net11 vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X31 gnd gnd vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X32 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X33 net4 net5 net5 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X34 net2 a_3720_130# net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X35 a_4940_2340# net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.25e+12p pd=1.2e+07u as=0p ps=0u w=1.5e+06u l=600000u
X36 net9 net9 net7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X37 gnd net10 net12 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X38 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X39 a_4500_160# v2 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X40 a_4940_160# gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=2.25e+12p pd=1.2e+07u as=0p ps=0u w=1.5e+06u l=600000u
X41 net1 net9 vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+12p ps=4e+07u w=1.5e+06u l=600000u
X42 net10 net9 a_4940_160# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X43 a_3720_130# a_3720_130# net4 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X44 net8 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X45 net6 v1 net11 vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X46 gnd net10 a_4940_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X47 vdd net9 a_4940_160# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X48 net16 gnd net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X49 net7 net5 net5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X50 gnd net9 net7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X51 net12 net10 gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X52 vout net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X53 net4 vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X54 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X55 net6 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X56 a_4060_800# gnd a_3720_130# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X57 a_4060_2340# vdd a_3720_130# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X58 vdd net10 net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X59 gnd net2 vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X60 net10 net10 net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X61 net13 vdd net6 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X62 a_4940_2340# net10 gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X63 net4 gnd a_4060_160# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X64 gnd gnd a_4500_160# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X65 vdd net9 net1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X66 gnd net9 net1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X67 net11 net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X68 vdd vdd net12 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X69 a_4940_160# net9 vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X70 vdd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X71 net6 vdd net22 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X72 vdd vdd gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X73 gnd gnd vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X74 net4 v2 net8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X75 net5 gnd net15 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X76 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X77 net9 vdd net10 vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X78 net2 vdd net13 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X79 gnd gnd vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X80 gnd net10 a_4940_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X81 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X82 net2 vout sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+07u
X83 vdd vdd a_4500_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X84 a_3720_130# a_3720_130# net7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X85 vout gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X86 net9 net10 a_4940_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X87 net7 v2 net11 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X88 a_4500_160# v1 net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X89 a_4500_2340# v1 net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X90 net1 net9 vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X91 a_4940_160# net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X92 net1 net9 net10 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X93 net3 net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X94 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X95 net12 net10 net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X96 vdd net9 a_4940_160# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X97 net3 net5 net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X98 net7 net9 net9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X99 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X100 a_4940_2340# vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X101 net8 gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X102 net15 gnd net3 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X103 net14 vdd net7 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X104 net10 vdd net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
.ends

*.subckt error_amp Cap1 Vref Vfb Cap2
X50k_res_0 VSUBS Vfb Cap1 k_res
Xopamp_0 Vref Vfb Cap2 opamp_0/vdd VSUBS opamp
*.ends

