*---------- DMG8601UFG Spice Model ----------
.SUBCKT power_nfet 10 20 30
*     TERMINALS:  D  G  S
M1 1 2 3 3  NMOS  L = 1 W = 1
RD 10 1 0.01441
RS 30 3 0.001
RG 20 2 202.6
CGS 2 3 1.466E-010
EGD 12 0 2 1 1
VFB 14 0 0
FFB 2 1  VFB 1
CGD 13 14 1E-009
R1 13 30 1
D1 12 13  DLIM
DDG 15 14  DCGD
R2 12 15 1
D2 15 0  DLIM
DSD 3 10  DSUB
.MODEL NMOS NMOS  LEVEL = 3  VMAX = 1.361E+005  ETA = 0.001  VTO = 0.8913
+ TOX = 6E-008  NSUB = 1E+016  KP = 97.33  KAPPA = 1  U0 = 400
.MODEL DCGD D  CJO = 2.802E-010  VJ = 0.2313  M = 0.4878
.MODEL DSUB D  IS = 2.098E-009  N = 1.133  RS = 0.02894  BV = 25  CJO = 2.541E-010  VJ = 0.1292  M = 0.32
.MODEL DLIM D  IS = 0.0001
.ENDS
