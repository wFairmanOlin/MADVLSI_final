magic
tech sky130A
timestamp 1620799792
<< nwell >>
rect 185 680 255 700
rect 185 615 255 635
rect 185 550 255 570
<< ndiff >>
rect 55 1085 80 1115
<< pdiffc >>
rect 185 680 255 700
rect 185 615 255 635
rect 185 550 255 570
<< poly >>
rect 0 5 40 15
rect 0 -10 10 5
rect -85 -15 10 -10
rect 30 -15 40 5
rect -85 -25 40 -15
rect -85 -170 2395 -160
rect -85 -175 2365 -170
rect 2355 -190 2365 -175
rect 2385 -190 2395 -170
rect 2355 -200 2395 -190
<< polycont >>
rect 10 -15 30 5
rect 2365 -190 2385 -170
<< locali >>
rect -85 1135 -55 1155
rect -80 1070 -55 1090
rect -80 625 -60 1070
rect -20 690 0 760
rect -80 -715 -55 625
rect -25 160 -5 625
rect 1020 270 1040 360
rect 2030 270 2050 360
rect 3040 270 3060 360
rect 4050 270 4070 360
rect -25 140 0 160
rect 0 5 40 15
rect 0 -15 10 5
rect 30 -5 40 5
rect 1975 -5 1995 145
rect 3050 140 3065 160
rect 30 -15 1995 -5
rect 0 -25 1995 -15
rect 2315 -110 2440 -75
rect 3035 -110 3055 140
rect 5080 75 5100 140
rect 5080 55 5135 75
rect 2355 -160 2375 -110
rect 2355 -170 2395 -160
rect 2355 -190 2365 -170
rect 2385 -190 2395 -170
rect 2355 -200 2395 -190
rect -80 -750 1525 -715
<< viali >>
rect 185 615 255 635
rect 5080 140 5100 160
<< metal1 >>
rect -80 580 75 625
rect -80 115 -40 580
rect 175 360 265 520
rect 5070 170 5115 175
rect 5070 135 5075 170
rect 5110 135 5115 170
rect 5070 130 5115 135
rect -80 15 10 115
<< via1 >>
rect 5075 160 5110 170
rect 5075 140 5080 160
rect 5080 140 5100 160
rect 5100 140 5110 160
rect 5075 135 5110 140
rect 1080 75 1115 110
<< metal2 >>
rect 5070 170 5115 175
rect 5070 135 5075 170
rect 5110 135 5115 170
rect 5070 130 5115 135
rect 1075 110 1120 115
rect 1075 75 1080 110
rect 1115 75 1120 110
rect 1075 70 1120 75
<< via2 >>
rect 5075 135 5110 170
rect 1080 75 1115 110
<< metal3 >>
rect 1165 115 1210 485
rect 5065 170 5115 180
rect 5065 135 5075 170
rect 5110 135 5115 170
rect 5065 125 5115 135
rect 1075 110 1210 115
rect 1075 75 1080 110
rect 1115 75 1210 110
rect 1075 70 1210 75
rect 1165 40 1210 70
<< via3 >>
rect 5075 135 5110 170
<< metal4 >>
rect 1090 435 5135 480
rect 5090 185 5135 435
rect 5075 175 5135 185
rect 5070 170 5135 175
rect 5070 135 5075 170
rect 5110 135 5135 170
rect 5070 130 5115 135
use 10k_res  10k_res_0
timestamp 1620799792
transform 0 1 2440 -1 0 -75
box 0 0 35 605
use and_gate_2p  and_gate_2p_0
timestamp 1620794368
transform 0 1 -155 -1 0 1050
box -275 100 535 445
use schmitt_inverter  schmitt_inverter_0 ~/Desktop
timestamp 1620698057
transform 1 0 120 0 1 15
box -120 -15 930 370
use schmitt_inverter  schmitt_inverter_1
timestamp 1620698057
transform 1 0 1130 0 1 15
box -120 -15 930 370
use schmitt_inverter  schmitt_inverter_2
timestamp 1620698057
transform 1 0 2140 0 1 15
box -120 -15 930 370
use schmitt_inverter  schmitt_inverter_3
timestamp 1620698057
transform 1 0 3150 0 1 15
box -120 -15 930 370
use schmitt_inverter  schmitt_inverter_4
timestamp 1620698057
transform 1 0 4160 0 1 15
box -120 -15 930 370
use 100k_res  100k_res_0
timestamp 1620671314
transform 0 1 1500 1 0 -615
box -135 25 540 815
use 4pf_cap  4pf_cap_0 ~/Desktop/MADVLSI_final/layout
timestamp 1620530160
transform 1 0 1315 0 1 1280
box -245 -800 3785 4275
<< labels >>
rlabel poly -85 -165 -85 -165 7 Cap2
port 1 w
rlabel poly -85 -20 -85 -20 7 Cap1
port 2 w
rlabel locali -85 1145 -85 1145 7 Enable
port 3 w
rlabel metal1 0 65 0 65 7 VN
port 4 w
rlabel metal1 175 445 175 445 7 VP
port 5 w
rlabel locali 5135 65 5135 65 3 Vclk
port 6 e
rlabel locali 3055 150 3055 150 7 net3
rlabel locali -80 1080 -80 1080 7 net4
rlabel locali -10 725 -10 725 1 net1
<< end >>
