magic
tech sky130A
timestamp 1620698057
<< nwell >>
rect -120 230 930 370
<< nmos >>
rect 130 0 145 100
rect 195 0 210 100
rect 260 0 275 100
rect 520 0 535 100
rect 585 0 600 100
rect 650 0 665 100
rect 715 0 730 100
<< pmos >>
rect 0 250 15 350
rect 65 250 80 350
rect 130 250 145 350
rect 195 250 210 350
rect 260 250 275 350
rect 325 250 340 350
rect 390 250 405 350
rect 455 250 470 350
rect 520 250 535 350
rect 585 250 600 350
rect 650 250 665 350
rect 715 250 730 350
rect 780 250 795 350
rect 845 250 860 350
<< ndiff >>
rect 80 85 130 100
rect 80 15 95 85
rect 115 15 130 85
rect 80 0 130 15
rect 145 85 195 100
rect 145 15 160 85
rect 180 15 195 85
rect 145 0 195 15
rect 210 85 260 100
rect 210 15 225 85
rect 245 15 260 85
rect 210 0 260 15
rect 275 85 325 100
rect 275 15 290 85
rect 310 15 325 85
rect 275 0 325 15
rect 470 85 520 100
rect 470 15 485 85
rect 505 15 520 85
rect 470 0 520 15
rect 535 85 585 100
rect 535 15 550 85
rect 570 15 585 85
rect 535 0 585 15
rect 600 85 650 100
rect 600 15 615 85
rect 635 15 650 85
rect 600 0 650 15
rect 665 85 715 100
rect 665 15 680 85
rect 700 15 715 85
rect 665 0 715 15
rect 730 85 780 100
rect 730 15 745 85
rect 765 15 780 85
rect 730 0 780 15
<< pdiff >>
rect -50 335 0 350
rect -50 265 -35 335
rect -15 265 0 335
rect -50 250 0 265
rect 15 335 65 350
rect 15 265 30 335
rect 50 265 65 335
rect 15 250 65 265
rect 80 335 130 350
rect 80 265 95 335
rect 115 265 130 335
rect 80 250 130 265
rect 145 335 195 350
rect 145 265 160 335
rect 180 265 195 335
rect 145 250 195 265
rect 210 335 260 350
rect 210 265 225 335
rect 245 265 260 335
rect 210 250 260 265
rect 275 335 325 350
rect 275 265 290 335
rect 310 265 325 335
rect 275 250 325 265
rect 340 335 390 350
rect 340 265 355 335
rect 375 265 390 335
rect 340 250 390 265
rect 405 335 455 350
rect 405 265 420 335
rect 440 265 455 335
rect 405 250 455 265
rect 470 335 520 350
rect 470 265 485 335
rect 505 265 520 335
rect 470 250 520 265
rect 535 335 585 350
rect 535 265 550 335
rect 570 265 585 335
rect 535 250 585 265
rect 600 335 650 350
rect 600 265 615 335
rect 635 265 650 335
rect 600 250 650 265
rect 665 335 715 350
rect 665 265 680 335
rect 700 265 715 335
rect 665 250 715 265
rect 730 335 780 350
rect 730 265 745 335
rect 765 265 780 335
rect 730 250 780 265
rect 795 335 845 350
rect 795 265 810 335
rect 830 265 845 335
rect 795 250 845 265
rect 860 335 910 350
rect 860 265 875 335
rect 895 265 910 335
rect 860 250 910 265
<< ndiffc >>
rect 95 15 115 85
rect 160 15 180 85
rect 225 15 245 85
rect 290 15 310 85
rect 485 15 505 85
rect 550 15 570 85
rect 615 15 635 85
rect 680 15 700 85
rect 745 15 765 85
<< pdiffc >>
rect -35 265 -15 335
rect 30 265 50 335
rect 95 265 115 335
rect 160 265 180 335
rect 225 265 245 335
rect 290 265 310 335
rect 355 265 375 335
rect 420 265 440 335
rect 485 265 505 335
rect 550 265 570 335
rect 615 265 635 335
rect 680 265 700 335
rect 745 265 765 335
rect 810 265 830 335
rect 875 265 895 335
<< psubdiff >>
rect 30 85 80 100
rect 30 15 45 85
rect 65 15 80 85
rect 30 0 80 15
rect 420 85 470 100
rect 420 15 435 85
rect 455 15 470 85
rect 420 0 470 15
<< nsubdiff >>
rect -100 335 -50 350
rect -100 265 -85 335
rect -65 265 -50 335
rect -100 250 -50 265
<< psubdiffcont >>
rect 45 15 65 85
rect 435 15 455 85
<< nsubdiffcont >>
rect -85 265 -65 335
<< poly >>
rect 0 350 15 365
rect 65 350 80 365
rect 130 350 145 365
rect 195 350 210 365
rect 260 350 275 365
rect 325 350 340 365
rect 390 350 405 365
rect 455 350 470 365
rect 520 350 535 365
rect 585 350 600 365
rect 650 350 665 365
rect 715 350 730 365
rect 780 350 795 365
rect 845 350 860 365
rect 0 235 15 250
rect 65 235 80 250
rect 130 235 145 250
rect 195 235 210 250
rect 0 220 210 235
rect -20 140 20 150
rect -20 120 -10 140
rect 10 125 20 140
rect 195 125 210 220
rect 10 120 210 125
rect -20 110 210 120
rect 130 100 145 110
rect 195 100 210 110
rect 260 235 275 250
rect 325 235 340 250
rect 260 220 340 235
rect 390 235 405 250
rect 455 235 470 250
rect 520 235 535 250
rect 585 235 600 250
rect 390 220 600 235
rect 260 100 275 220
rect 325 210 365 220
rect 325 190 335 210
rect 355 190 365 210
rect 325 180 365 190
rect 390 155 405 220
rect 300 145 405 155
rect 300 125 310 145
rect 330 140 405 145
rect 330 125 340 140
rect 585 125 600 220
rect 650 235 665 250
rect 715 235 730 250
rect 780 235 795 250
rect 845 235 860 250
rect 650 220 860 235
rect 650 165 665 220
rect 625 155 665 165
rect 625 135 635 155
rect 655 135 665 155
rect 625 125 665 135
rect 300 115 340 125
rect 520 110 600 125
rect 520 100 535 110
rect 585 100 600 110
rect 650 110 730 125
rect 650 100 665 110
rect 715 100 730 110
rect 130 -15 145 0
rect 195 -15 210 0
rect 260 -15 275 0
rect 520 -15 535 0
rect 585 -15 600 0
rect 650 -15 665 0
rect 715 -15 730 0
<< polycont >>
rect -10 120 10 140
rect 335 190 355 210
rect 310 125 330 145
rect 635 135 655 155
<< locali >>
rect -95 335 -5 345
rect -95 265 -85 335
rect -65 265 -35 335
rect -15 265 -5 335
rect -95 255 -5 265
rect 20 335 60 345
rect 20 265 30 335
rect 50 265 60 335
rect 20 255 60 265
rect 85 335 125 345
rect 85 265 95 335
rect 115 265 125 335
rect 85 255 125 265
rect 150 335 190 345
rect 150 265 160 335
rect 180 265 190 335
rect 150 255 190 265
rect 215 335 255 345
rect 215 265 225 335
rect 245 265 255 335
rect 215 255 255 265
rect 280 335 320 345
rect 280 265 290 335
rect 310 265 320 335
rect 280 255 320 265
rect 345 335 385 345
rect 345 265 355 335
rect 375 265 385 335
rect 345 255 385 265
rect 410 335 450 345
rect 410 265 420 335
rect 440 265 450 335
rect 410 255 450 265
rect 475 335 515 345
rect 475 265 485 335
rect 505 265 515 335
rect 475 255 515 265
rect 540 335 580 345
rect 540 265 550 335
rect 570 265 580 335
rect 540 255 580 265
rect 605 335 645 345
rect 605 265 615 335
rect 635 265 645 335
rect 605 255 645 265
rect 670 335 710 345
rect 670 265 680 335
rect 700 265 710 335
rect 670 255 710 265
rect 735 335 775 345
rect 735 265 745 335
rect 765 265 775 335
rect 735 255 775 265
rect 800 335 840 345
rect 800 265 810 335
rect 830 265 840 335
rect 800 255 840 265
rect 865 335 905 345
rect 865 265 875 335
rect 895 265 905 335
rect 865 255 905 265
rect 40 235 60 255
rect 150 235 170 255
rect 40 215 170 235
rect 150 155 170 215
rect 280 155 300 255
rect 430 235 450 255
rect 540 235 560 255
rect 325 210 365 220
rect 430 215 560 235
rect 325 190 335 210
rect 355 200 365 210
rect 355 195 405 200
rect 540 195 560 215
rect 355 190 560 195
rect 325 180 560 190
rect 365 175 560 180
rect -20 145 20 150
rect -120 140 20 145
rect -120 125 -10 140
rect -20 120 -10 125
rect 10 120 20 140
rect -20 110 20 120
rect 150 145 340 155
rect 150 135 310 145
rect 150 95 170 135
rect 280 125 310 135
rect 330 125 340 145
rect 280 115 340 125
rect 540 145 560 175
rect 690 235 710 255
rect 800 235 820 255
rect 690 215 820 235
rect 625 155 665 165
rect 625 145 635 155
rect 540 135 635 145
rect 655 135 665 155
rect 540 125 665 135
rect 690 145 710 215
rect 690 125 930 145
rect 280 95 300 115
rect 540 95 560 125
rect 690 95 710 125
rect 35 85 125 95
rect 35 15 45 85
rect 65 15 95 85
rect 115 15 125 85
rect 35 5 125 15
rect 150 85 190 95
rect 150 15 160 85
rect 180 15 190 85
rect 150 5 190 15
rect 215 85 255 95
rect 215 15 225 85
rect 245 15 255 85
rect 215 5 255 15
rect 280 85 320 95
rect 280 15 290 85
rect 310 15 320 85
rect 280 5 320 15
rect 425 85 515 95
rect 425 15 435 85
rect 455 15 485 85
rect 505 15 515 85
rect 425 5 515 15
rect 540 85 580 95
rect 540 15 550 85
rect 570 15 580 85
rect 540 5 580 15
rect 605 85 645 95
rect 605 15 615 85
rect 635 15 645 85
rect 605 5 645 15
rect 670 85 710 95
rect 670 15 680 85
rect 700 15 710 85
rect 670 5 710 15
rect 735 85 775 95
rect 735 15 745 85
rect 765 15 775 85
rect 735 5 775 15
<< viali >>
rect -85 265 -65 335
rect -35 265 -15 335
rect 95 265 115 335
rect 225 265 245 335
rect 355 265 375 335
rect 485 265 505 335
rect 615 265 635 335
rect 745 265 765 335
rect 875 265 895 335
rect 45 15 65 85
rect 95 15 115 85
rect 225 15 245 85
rect 435 15 455 85
rect 485 15 505 85
rect 615 15 635 85
rect 745 15 765 85
<< metal1 >>
rect -120 335 930 350
rect -120 265 -85 335
rect -65 265 -35 335
rect -15 265 95 335
rect 115 265 225 335
rect 245 265 355 335
rect 375 265 485 335
rect 505 265 615 335
rect 635 265 745 335
rect 765 265 875 335
rect 895 265 930 335
rect -120 250 930 265
rect -120 85 930 100
rect -120 15 45 85
rect 65 15 95 85
rect 115 15 225 85
rect 245 15 435 85
rect 455 15 485 85
rect 505 15 615 85
rect 635 15 745 85
rect 765 15 930 85
rect -120 0 930 15
<< labels >>
rlabel metal1 -120 50 -120 50 7 VN
port 4 w
rlabel metal1 -120 295 -120 295 7 VP
port 3 w
rlabel locali 930 135 930 135 3 Z
port 2 e
rlabel locali -120 135 -120 135 7 A
port 1 w
<< end >>
