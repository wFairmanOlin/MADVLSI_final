*SRC=DMN3150LW;DI_DMN3150LW;MOSFETs N;Enh;28.0V 1.60A 88.0mohms  Diodes Inc MOSFET
*SYM=POWMOSN
.SUBCKT power_nfet   10 20 30
*     TERMINALS:  D  G  S
M1   1  2  3  3  DMOS L=1 W=1
RD  10  1  40.8m
RS  40  3  3.20m
RG  20  2  93.7
CGS  2  3  257p
EGD 12  0  2  1  1
VFB 14  0  0
FFB  2  1  VFB  1
CGD 13 14  219p
R1  13  0  1.00
D1  12 13  DLIM
DDG 15 14  DCGD
R2  12 15  1.00
D2  15  0  DLIM
DSD  3 10  DSUB
LS  30 40  7.50n
.MODEL DMOS NMOS(LEVEL=3 VMAX=58.3k THETA=80.0m
+ ETA=2.00m VTO=1.40 KP=21.8
.MODEL DCGD D (CJO=219p VJ=0.600 M=0.680
.MODEL DSUB D (IS=6.64n N=1.50 RS=0.256 BV=28.0
+ CJO=85.0p VJ=0.800 M=0.420 TT=162n
.MODEL DLIM D (IS=100U)
.ends
