magic
tech sky130A
timestamp 1620808523
<< locali >>
rect -50 725 -10 1315
rect -50 705 -40 725
rect -20 705 -10 725
rect -50 695 -10 705
rect -725 -10 -690 0
<< viali >>
rect -40 705 -20 725
<< metal1 >>
rect -50 725 30 735
rect -50 705 -40 725
rect -20 705 30 725
rect -50 695 30 705
rect 5640 395 5655 435
rect 5640 305 5655 345
rect 5640 245 5655 285
use 250k_res  250k_res_0
timestamp 1620673804
transform 1 0 -725 0 1 0
box 0 0 675 1315
use opamp  opamp_0 ~/Desktop/MADVLSI_final/layout
timestamp 1620660520
transform 1 0 230 0 1 -30
box -230 30 5425 1700
<< labels >>
rlabel locali -710 -10 -710 -10 1 Cap1
port 1 n
rlabel metal1 5655 325 5655 325 3 Vref
port 2 e
rlabel metal1 5640 245 5655 285 3 Vfb
port 3 e
rlabel metal1 5655 415 5655 415 3 Cap2
port 4 e
<< end >>
