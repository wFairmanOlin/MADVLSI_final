* SPICE3 file created from opamp_square.ext - technology: sky130A

X0 gnd gnd vout gnd sky130_fd_pr__nfet_01v8 ad=1.2e+13p pd=6.4e+07u as=3e+12p ps=1.6e+07u w=1.5e+06u l=600000u
X1 net16 gnd net4 gnd sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=4e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X2 a_3720_110# a_3720_110# net7 gnd sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=4e+06u as=3e+12p ps=1.6e+07u w=1.5e+06u l=600000u
X3 net2 a_3720_110# net3 vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X4 vout net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X5 net6 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X6 net7 vdd a_4060_2340# vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X7 vdd net10 net12 vdd sky130_fd_pr__pfet_01v8 ad=1.2e+13p pd=6.4e+07u as=2.25e+12p ps=1.2e+07u w=1.5e+06u l=600000u
X8 vdd vdd net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=3e+12p ps=1.6e+07u w=1.5e+06u l=600000u
X9 a_4500_140# v1 net3 gnd sky130_fd_pr__nfet_01v8 ad=1.5e+12p pd=8e+06u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X10 gnd net2 vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X11 a_4940_140# net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=2.25e+12p pd=1.2e+07u as=0p ps=0u w=1.5e+06u l=600000u
X12 net1 net9 net10 gnd sky130_fd_pr__nfet_01v8 ad=2.25e+12p pd=1.2e+07u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X13 net4 gnd a_4060_140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X14 net4 net10 net10 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X15 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=3e+12p pd=1.6e+07u as=0p ps=0u w=1.5e+06u l=600000u
X16 net5 vdd net14 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X17 gnd gnd a_4500_140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X18 vdd net9 net1 gnd sky130_fd_pr__nfet_01v8 ad=7.5e+12p pd=4e+07u as=0p ps=0u w=1.5e+06u l=600000u
X19 vdd net10 a_4500_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X20 gnd vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=7.5e+12p pd=4e+07u as=0p ps=0u w=1.5e+06u l=600000u
X21 net7 net9 net9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X22 net22 vdd net2 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X23 net15 gnd net3 gnd sky130_fd_pr__nfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X24 net12 net10 gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X25 vdd net10 net3 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X26 a_4940_140# net9 vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X27 vdd gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X28 gnd gnd vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X29 a_4500_2340# v2 net7 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X30 vout net2 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X31 net4 net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X32 net4 v2 net8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X33 net7 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X34 gnd net2 vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X35 net11 vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X36 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X37 net4 net5 net5 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X38 net3 gnd a_4060_780# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X39 a_4940_2340# net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=2.25e+12p pd=1.2e+07u as=0p ps=0u w=1.5e+06u l=600000u
X40 vout gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X41 gnd net9 a_4500_140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X42 net10 gnd net9 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X43 gnd net10 net12 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X44 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X45 net1 net9 vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X46 net7 gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X47 net9 gnd net10 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X48 a_3720_110# a_3720_110# net4 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X49 gnd gnd net7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X50 net3 v1 net8 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X51 net6 v1 net11 vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X52 vdd net9 a_4940_140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X53 gnd net10 a_4940_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X54 net8 gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X55 net2 vout sky130_fd_pr__cap_mim_m3_1 l=1.2e+07u w=2e+07u
X56 vout gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X57 net12 net10 gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X58 net4 vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X59 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X60 net6 net5 net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=1.5e+12p ps=8e+06u w=1.5e+06u l=600000u
X61 a_4060_2340# vdd a_3720_110# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X62 gnd net9 net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X63 net9 net9 net7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X64 vdd net10 net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X65 net10 net10 net4 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X66 a_4060_140# gnd net2 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X67 net13 vdd net6 vdd sky130_fd_pr__pfet_01v8 ad=7.5e+11p pd=4e+06u as=0p ps=0u w=1.5e+06u l=600000u
X68 a_4940_2340# net10 gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X69 net10 net9 a_4940_140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X70 net11 net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X71 net8 net9 gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X72 gnd gnd net1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X73 vdd vdd net12 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X74 net6 vdd net22 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X75 vdd vdd gnd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X76 net7 net5 net5 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=7.5e+11p ps=4e+06u w=1.5e+06u l=600000u
X77 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X78 net9 vdd net10 vdd sky130_fd_pr__pfet_01v8 ad=1.5e+12p pd=8e+06u as=0p ps=0u w=1.5e+06u l=600000u
X79 gnd net9 net7 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X80 net2 vdd net13 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X81 gnd net10 a_4940_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X82 vout net2 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X83 net2 gnd net16 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X84 a_4060_780# gnd a_3720_110# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X85 vdd vdd a_4500_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X86 gnd gnd vout gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X87 net9 net10 a_4940_2340# vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X88 net7 v2 net11 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X89 net2 a_3720_110# net6 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X90 a_4500_2340# v1 net6 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X91 gnd net9 net1 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X92 net3 net10 vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X93 a_4500_140# v2 net4 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X94 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X95 net12 net10 net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X96 a_4940_140# gnd gnd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X97 net1 net9 vdd gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X98 net3 net5 net2 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X99 vdd net2 vout vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X100 a_4940_2340# vdd vdd vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X101 net5 gnd net15 gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X102 vdd net9 a_4940_140# gnd sky130_fd_pr__nfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X103 net14 vdd net7 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u
X104 net10 vdd net9 vdd sky130_fd_pr__pfet_01v8 ad=0p pd=0u as=0p ps=0u w=1.5e+06u l=600000u

