.subckt sky130_fd_pr__pnp_05v0  E B C
*.iopin E
*.iopin B
*.iopin C
XQ1 C B E C sky130_fd_pr__pnp_05v5_W0p68L0p68
.ends
