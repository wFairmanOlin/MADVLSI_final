magic
tech sky130A
magscale 1 2
timestamp 1620823543
<< nwell >>
rect 7280 1950 8040 6350
<< pwell >>
rect -1110 -637 -334 -484
rect -1110 -1127 -977 -637
rect -487 -1127 -334 -637
rect -1110 -1280 -334 -1127
rect -310 -637 486 -484
rect -310 -1127 -157 -637
rect 333 -1127 486 -637
rect -310 -1280 486 -1127
rect 510 -637 1306 -484
rect 510 -1127 663 -637
rect 1153 -1127 1306 -637
rect 510 -1280 1306 -1127
rect 1330 -637 2126 -484
rect 1330 -1127 1483 -637
rect 1973 -1127 2126 -637
rect 1330 -1280 2126 -1127
rect 2150 -637 2946 -484
rect 2150 -1127 2303 -637
rect 2793 -1127 2946 -637
rect 2150 -1280 2946 -1127
rect 2970 -637 3766 -484
rect 2970 -1127 3123 -637
rect 3613 -1127 3766 -637
rect 2970 -1280 3766 -1127
rect 3790 -637 4586 -484
rect 3790 -1127 3943 -637
rect 4433 -1127 4586 -637
rect 3790 -1280 4586 -1127
rect 4610 -637 5406 -484
rect 4610 -1127 4763 -637
rect 5253 -1127 5406 -637
rect 4610 -1280 5406 -1127
rect 5430 -637 6226 -484
rect 5430 -1127 5583 -637
rect 6073 -1127 6226 -637
rect 5430 -1280 6226 -1127
rect 6250 -637 7046 -484
rect 6250 -1127 6403 -637
rect 6893 -1127 7046 -637
rect 6250 -1280 7046 -1127
rect 7100 -637 7896 -484
rect 7100 -1127 7253 -637
rect 7743 -1127 7896 -637
rect 7100 -1280 7896 -1127
rect -1110 -1457 -334 -1304
rect -1110 -1947 -977 -1457
rect -487 -1947 -334 -1457
rect -1110 -2100 -334 -1947
rect -310 -1457 486 -1304
rect -310 -1947 -157 -1457
rect 333 -1947 486 -1457
rect -310 -2100 486 -1947
rect 510 -1457 1306 -1304
rect 510 -1947 663 -1457
rect 1153 -1947 1306 -1457
rect 510 -2100 1306 -1947
rect 1330 -1457 2126 -1304
rect 1330 -1947 1483 -1457
rect 1973 -1947 2126 -1457
rect 1330 -2100 2126 -1947
rect 2150 -1457 2946 -1304
rect 2150 -1947 2303 -1457
rect 2793 -1947 2946 -1457
rect 2150 -2100 2946 -1947
rect 2970 -1457 3766 -1304
rect 2970 -1947 3123 -1457
rect 3613 -1947 3766 -1457
rect 2970 -2100 3766 -1947
rect 3790 -1457 4586 -1304
rect 3790 -1947 3943 -1457
rect 4433 -1947 4586 -1457
rect 3790 -2100 4586 -1947
rect 4610 -1457 5406 -1304
rect 4610 -1947 4763 -1457
rect 5253 -1947 5406 -1457
rect 4610 -2100 5406 -1947
rect 5430 -1457 6226 -1304
rect 5430 -1947 5583 -1457
rect 6073 -1947 6226 -1457
rect 5430 -2100 6226 -1947
rect 6250 -1457 7046 -1304
rect 6250 -1947 6403 -1457
rect 6893 -1947 7046 -1457
rect 6250 -2100 7046 -1947
rect -1110 -2277 -334 -2124
rect -1110 -2767 -977 -2277
rect -487 -2767 -334 -2277
rect -1110 -2920 -334 -2767
rect -310 -2277 486 -2124
rect -310 -2767 -157 -2277
rect 333 -2767 486 -2277
rect -310 -2920 486 -2767
rect 510 -2277 1306 -2124
rect 510 -2767 663 -2277
rect 1153 -2767 1306 -2277
rect 510 -2920 1306 -2767
rect 1330 -2277 2126 -2124
rect 1330 -2767 1483 -2277
rect 1973 -2767 2126 -2277
rect 1330 -2920 2126 -2767
rect 2150 -2277 2946 -2124
rect 2150 -2767 2303 -2277
rect 2793 -2767 2946 -2277
rect 2150 -2920 2946 -2767
rect 2970 -2277 3766 -2124
rect 2970 -2767 3123 -2277
rect 3613 -2767 3766 -2277
rect 2970 -2920 3766 -2767
rect 3790 -2277 4586 -2124
rect 3790 -2767 3943 -2277
rect 4433 -2767 4586 -2277
rect 3790 -2920 4586 -2767
rect 4610 -2277 5406 -2124
rect 4610 -2767 4763 -2277
rect 5253 -2767 5406 -2277
rect 4610 -2920 5406 -2767
rect 5430 -2277 6226 -2124
rect 5430 -2767 5583 -2277
rect 6073 -2767 6226 -2277
rect 5430 -2920 6226 -2767
rect 6250 -2277 7046 -2124
rect 6250 -2767 6403 -2277
rect 6893 -2767 7046 -2277
rect 6250 -2920 7046 -2767
rect -1110 -3097 -334 -2944
rect -1110 -3587 -977 -3097
rect -487 -3587 -334 -3097
rect -1110 -3740 -334 -3587
rect -310 -3097 486 -2944
rect -310 -3587 -157 -3097
rect 333 -3587 486 -3097
rect -310 -3740 486 -3587
rect 510 -3097 1306 -2944
rect 510 -3587 663 -3097
rect 1153 -3587 1306 -3097
rect 510 -3740 1306 -3587
rect 1330 -3097 2126 -2944
rect 1330 -3587 1483 -3097
rect 1973 -3587 2126 -3097
rect 1330 -3740 2126 -3587
rect 2150 -3097 2946 -2944
rect 2150 -3587 2303 -3097
rect 2793 -3587 2946 -3097
rect 2150 -3740 2946 -3587
rect 2970 -3097 3766 -2944
rect 2970 -3587 3123 -3097
rect 3613 -3587 3766 -3097
rect 2970 -3740 3766 -3587
rect 3790 -3097 4586 -2944
rect 3790 -3587 3943 -3097
rect 4433 -3587 4586 -3097
rect 3790 -3740 4586 -3587
rect 4610 -3097 5406 -2944
rect 4610 -3587 4763 -3097
rect 5253 -3587 5406 -3097
rect 4610 -3740 5406 -3587
rect 5430 -3097 6226 -2944
rect 5430 -3587 5583 -3097
rect 6073 -3587 6226 -3097
rect 5430 -3740 6226 -3587
rect 6250 -3097 7046 -2944
rect 6250 -3587 6403 -3097
rect 6893 -3587 7046 -3097
rect 6250 -3740 7046 -3587
rect -1110 -3917 -334 -3764
rect -1110 -4407 -977 -3917
rect -487 -4407 -334 -3917
rect -1110 -4560 -334 -4407
rect -310 -3917 486 -3764
rect -310 -4407 -157 -3917
rect 333 -4407 486 -3917
rect -310 -4560 486 -4407
rect 510 -3917 1306 -3764
rect 510 -4407 663 -3917
rect 1153 -4407 1306 -3917
rect 510 -4560 1306 -4407
rect 1330 -3917 2126 -3764
rect 1330 -4407 1483 -3917
rect 1973 -4407 2126 -3917
rect 1330 -4560 2126 -4407
rect 2150 -3917 2946 -3764
rect 2150 -4407 2303 -3917
rect 2793 -4407 2946 -3917
rect 2150 -4560 2946 -4407
rect 2970 -3917 3766 -3764
rect 2970 -4407 3123 -3917
rect 3613 -4407 3766 -3917
rect 2970 -4560 3766 -4407
rect 3790 -3917 4586 -3764
rect 3790 -4407 3943 -3917
rect 4433 -4407 4586 -3917
rect 3790 -4560 4586 -4407
rect 4610 -3917 5406 -3764
rect 4610 -4407 4763 -3917
rect 5253 -4407 5406 -3917
rect 4610 -4560 5406 -4407
rect 5430 -3917 6226 -3764
rect 5430 -4407 5583 -3917
rect 6073 -4407 6226 -3917
rect 5430 -4560 6226 -4407
rect 6250 -3917 7046 -3764
rect 6250 -4407 6403 -3917
rect 6893 -4407 7046 -3917
rect 6250 -4560 7046 -4407
<< nbase >>
rect -977 -1127 -487 -637
rect -157 -1127 333 -637
rect 663 -1127 1153 -637
rect 1483 -1127 1973 -637
rect 2303 -1127 2793 -637
rect 3123 -1127 3613 -637
rect 3943 -1127 4433 -637
rect 4763 -1127 5253 -637
rect 5583 -1127 6073 -637
rect 6403 -1127 6893 -637
rect 7253 -1127 7743 -637
rect -977 -1947 -487 -1457
rect -157 -1947 333 -1457
rect 663 -1947 1153 -1457
rect 1483 -1947 1973 -1457
rect 2303 -1947 2793 -1457
rect 3123 -1947 3613 -1457
rect 3943 -1947 4433 -1457
rect 4763 -1947 5253 -1457
rect 5583 -1947 6073 -1457
rect 6403 -1947 6893 -1457
rect -977 -2767 -487 -2277
rect -157 -2767 333 -2277
rect 663 -2767 1153 -2277
rect 1483 -2767 1973 -2277
rect 2303 -2767 2793 -2277
rect 3123 -2767 3613 -2277
rect 3943 -2767 4433 -2277
rect 4763 -2767 5253 -2277
rect 5583 -2767 6073 -2277
rect 6403 -2767 6893 -2277
rect -977 -3587 -487 -3097
rect -157 -3587 333 -3097
rect 663 -3587 1153 -3097
rect 1483 -3587 1973 -3097
rect 2303 -3587 2793 -3097
rect 3123 -3587 3613 -3097
rect 3943 -3587 4433 -3097
rect 4763 -3587 5253 -3097
rect 5583 -3587 6073 -3097
rect 6403 -3587 6893 -3097
rect -977 -4407 -487 -3917
rect -157 -4407 333 -3917
rect 663 -4407 1153 -3917
rect 1483 -4407 1973 -3917
rect 2303 -4407 2793 -3917
rect 3123 -4407 3613 -3917
rect 3943 -4407 4433 -3917
rect 4763 -4407 5253 -3917
rect 5583 -4407 6073 -3917
rect 6403 -4407 6893 -3917
<< pmos >>
rect 7500 4270 7530 6270
rect 7830 4270 7860 6270
rect 7500 2060 7530 4060
rect 7830 2060 7860 4060
<< pdiff >>
rect 7400 6240 7500 6270
rect 7400 4300 7430 6240
rect 7470 4300 7500 6240
rect 7400 4270 7500 4300
rect 7530 6240 7630 6270
rect 7730 6240 7830 6270
rect 7530 4300 7560 6240
rect 7600 4300 7630 6240
rect 7730 4300 7760 6240
rect 7800 4300 7830 6240
rect 7530 4270 7630 4300
rect 7730 4270 7830 4300
rect 7860 6240 7960 6270
rect 7860 4300 7890 6240
rect 7930 4300 7960 6240
rect 7860 4270 7960 4300
rect 7400 4030 7500 4060
rect 7400 2090 7430 4030
rect 7470 2090 7500 4030
rect 7400 2060 7500 2090
rect 7530 4030 7630 4060
rect 7730 4030 7830 4060
rect 7530 2090 7560 4030
rect 7600 2090 7630 4030
rect 7730 2090 7760 4030
rect 7800 2090 7830 4030
rect 7530 2060 7630 2090
rect 7730 2060 7830 2090
rect 7860 4030 7960 4060
rect 7860 2090 7890 4030
rect 7930 2090 7960 4030
rect 7860 2060 7960 2090
rect -800 -831 -664 -814
rect -800 -933 -783 -831
rect -681 -933 -664 -831
rect -800 -950 -664 -933
rect 20 -831 156 -814
rect 20 -933 37 -831
rect 139 -933 156 -831
rect 20 -950 156 -933
rect 840 -831 976 -814
rect 840 -933 857 -831
rect 959 -933 976 -831
rect 840 -950 976 -933
rect 1660 -831 1796 -814
rect 1660 -933 1677 -831
rect 1779 -933 1796 -831
rect 1660 -950 1796 -933
rect 2480 -831 2616 -814
rect 2480 -933 2497 -831
rect 2599 -933 2616 -831
rect 2480 -950 2616 -933
rect 3300 -831 3436 -814
rect 3300 -933 3317 -831
rect 3419 -933 3436 -831
rect 3300 -950 3436 -933
rect 4120 -831 4256 -814
rect 4120 -933 4137 -831
rect 4239 -933 4256 -831
rect 4120 -950 4256 -933
rect 4940 -831 5076 -814
rect 4940 -933 4957 -831
rect 5059 -933 5076 -831
rect 4940 -950 5076 -933
rect 5760 -831 5896 -814
rect 5760 -933 5777 -831
rect 5879 -933 5896 -831
rect 5760 -950 5896 -933
rect 6580 -831 6716 -814
rect 6580 -933 6597 -831
rect 6699 -933 6716 -831
rect 6580 -950 6716 -933
rect 7430 -831 7566 -814
rect 7430 -933 7447 -831
rect 7549 -933 7566 -831
rect 7430 -950 7566 -933
rect -800 -1651 -664 -1634
rect -800 -1753 -783 -1651
rect -681 -1753 -664 -1651
rect -800 -1770 -664 -1753
rect 20 -1651 156 -1634
rect 20 -1753 37 -1651
rect 139 -1753 156 -1651
rect 20 -1770 156 -1753
rect 840 -1651 976 -1634
rect 840 -1753 857 -1651
rect 959 -1753 976 -1651
rect 840 -1770 976 -1753
rect 1660 -1651 1796 -1634
rect 1660 -1753 1677 -1651
rect 1779 -1753 1796 -1651
rect 1660 -1770 1796 -1753
rect 2480 -1651 2616 -1634
rect 2480 -1753 2497 -1651
rect 2599 -1753 2616 -1651
rect 2480 -1770 2616 -1753
rect 3300 -1651 3436 -1634
rect 3300 -1753 3317 -1651
rect 3419 -1753 3436 -1651
rect 3300 -1770 3436 -1753
rect 4120 -1651 4256 -1634
rect 4120 -1753 4137 -1651
rect 4239 -1753 4256 -1651
rect 4120 -1770 4256 -1753
rect 4940 -1651 5076 -1634
rect 4940 -1753 4957 -1651
rect 5059 -1753 5076 -1651
rect 4940 -1770 5076 -1753
rect 5760 -1651 5896 -1634
rect 5760 -1753 5777 -1651
rect 5879 -1753 5896 -1651
rect 5760 -1770 5896 -1753
rect 6580 -1651 6716 -1634
rect 6580 -1753 6597 -1651
rect 6699 -1753 6716 -1651
rect 6580 -1770 6716 -1753
rect -800 -2471 -664 -2454
rect -800 -2573 -783 -2471
rect -681 -2573 -664 -2471
rect -800 -2590 -664 -2573
rect 20 -2471 156 -2454
rect 20 -2573 37 -2471
rect 139 -2573 156 -2471
rect 20 -2590 156 -2573
rect 840 -2471 976 -2454
rect 840 -2573 857 -2471
rect 959 -2573 976 -2471
rect 840 -2590 976 -2573
rect 1660 -2471 1796 -2454
rect 1660 -2573 1677 -2471
rect 1779 -2573 1796 -2471
rect 1660 -2590 1796 -2573
rect 2480 -2471 2616 -2454
rect 2480 -2573 2497 -2471
rect 2599 -2573 2616 -2471
rect 2480 -2590 2616 -2573
rect 3300 -2471 3436 -2454
rect 3300 -2573 3317 -2471
rect 3419 -2573 3436 -2471
rect 3300 -2590 3436 -2573
rect 4120 -2471 4256 -2454
rect 4120 -2573 4137 -2471
rect 4239 -2573 4256 -2471
rect 4120 -2590 4256 -2573
rect 4940 -2471 5076 -2454
rect 4940 -2573 4957 -2471
rect 5059 -2573 5076 -2471
rect 4940 -2590 5076 -2573
rect 5760 -2471 5896 -2454
rect 5760 -2573 5777 -2471
rect 5879 -2573 5896 -2471
rect 5760 -2590 5896 -2573
rect 6580 -2471 6716 -2454
rect 6580 -2573 6597 -2471
rect 6699 -2573 6716 -2471
rect 6580 -2590 6716 -2573
rect -800 -3291 -664 -3274
rect -800 -3393 -783 -3291
rect -681 -3393 -664 -3291
rect -800 -3410 -664 -3393
rect 20 -3291 156 -3274
rect 20 -3393 37 -3291
rect 139 -3393 156 -3291
rect 20 -3410 156 -3393
rect 840 -3291 976 -3274
rect 840 -3393 857 -3291
rect 959 -3393 976 -3291
rect 840 -3410 976 -3393
rect 1660 -3291 1796 -3274
rect 1660 -3393 1677 -3291
rect 1779 -3393 1796 -3291
rect 1660 -3410 1796 -3393
rect 2480 -3291 2616 -3274
rect 2480 -3393 2497 -3291
rect 2599 -3393 2616 -3291
rect 2480 -3410 2616 -3393
rect 3300 -3291 3436 -3274
rect 3300 -3393 3317 -3291
rect 3419 -3393 3436 -3291
rect 3300 -3410 3436 -3393
rect 4120 -3291 4256 -3274
rect 4120 -3393 4137 -3291
rect 4239 -3393 4256 -3291
rect 4120 -3410 4256 -3393
rect 4940 -3291 5076 -3274
rect 4940 -3393 4957 -3291
rect 5059 -3393 5076 -3291
rect 4940 -3410 5076 -3393
rect 5760 -3291 5896 -3274
rect 5760 -3393 5777 -3291
rect 5879 -3393 5896 -3291
rect 5760 -3410 5896 -3393
rect 6580 -3291 6716 -3274
rect 6580 -3393 6597 -3291
rect 6699 -3393 6716 -3291
rect 6580 -3410 6716 -3393
rect -800 -4111 -664 -4094
rect -800 -4213 -783 -4111
rect -681 -4213 -664 -4111
rect -800 -4230 -664 -4213
rect 20 -4111 156 -4094
rect 20 -4213 37 -4111
rect 139 -4213 156 -4111
rect 20 -4230 156 -4213
rect 840 -4111 976 -4094
rect 840 -4213 857 -4111
rect 959 -4213 976 -4111
rect 840 -4230 976 -4213
rect 1660 -4111 1796 -4094
rect 1660 -4213 1677 -4111
rect 1779 -4213 1796 -4111
rect 1660 -4230 1796 -4213
rect 2480 -4111 2616 -4094
rect 2480 -4213 2497 -4111
rect 2599 -4213 2616 -4111
rect 2480 -4230 2616 -4213
rect 3300 -4111 3436 -4094
rect 3300 -4213 3317 -4111
rect 3419 -4213 3436 -4111
rect 3300 -4230 3436 -4213
rect 4120 -4111 4256 -4094
rect 4120 -4213 4137 -4111
rect 4239 -4213 4256 -4111
rect 4120 -4230 4256 -4213
rect 4940 -4111 5076 -4094
rect 4940 -4213 4957 -4111
rect 5059 -4213 5076 -4111
rect 4940 -4230 5076 -4213
rect 5760 -4111 5896 -4094
rect 5760 -4213 5777 -4111
rect 5879 -4213 5896 -4111
rect 5760 -4230 5896 -4213
rect 6580 -4111 6716 -4094
rect 6580 -4213 6597 -4111
rect 6699 -4213 6716 -4111
rect 6580 -4230 6716 -4213
<< pdiffc >>
rect 7430 4300 7470 6240
rect 7560 4300 7600 6240
rect 7760 4300 7800 6240
rect 7890 4300 7930 6240
rect 7430 2090 7470 4030
rect 7560 2090 7600 4030
rect 7760 2090 7800 4030
rect 7890 2090 7930 4030
rect -783 -933 -681 -831
rect 37 -933 139 -831
rect 857 -933 959 -831
rect 1677 -933 1779 -831
rect 2497 -933 2599 -831
rect 3317 -933 3419 -831
rect 4137 -933 4239 -831
rect 4957 -933 5059 -831
rect 5777 -933 5879 -831
rect 6597 -933 6699 -831
rect 7447 -933 7549 -831
rect -783 -1753 -681 -1651
rect 37 -1753 139 -1651
rect 857 -1753 959 -1651
rect 1677 -1753 1779 -1651
rect 2497 -1753 2599 -1651
rect 3317 -1753 3419 -1651
rect 4137 -1753 4239 -1651
rect 4957 -1753 5059 -1651
rect 5777 -1753 5879 -1651
rect 6597 -1753 6699 -1651
rect -783 -2573 -681 -2471
rect 37 -2573 139 -2471
rect 857 -2573 959 -2471
rect 1677 -2573 1779 -2471
rect 2497 -2573 2599 -2471
rect 3317 -2573 3419 -2471
rect 4137 -2573 4239 -2471
rect 4957 -2573 5059 -2471
rect 5777 -2573 5879 -2471
rect 6597 -2573 6699 -2471
rect -783 -3393 -681 -3291
rect 37 -3393 139 -3291
rect 857 -3393 959 -3291
rect 1677 -3393 1779 -3291
rect 2497 -3393 2599 -3291
rect 3317 -3393 3419 -3291
rect 4137 -3393 4239 -3291
rect 4957 -3393 5059 -3291
rect 5777 -3393 5879 -3291
rect 6597 -3393 6699 -3291
rect -783 -4213 -681 -4111
rect 37 -4213 139 -4111
rect 857 -4213 959 -4111
rect 1677 -4213 1779 -4111
rect 2497 -4213 2599 -4111
rect 3317 -4213 3419 -4111
rect 4137 -4213 4239 -4111
rect 4957 -4213 5059 -4111
rect 5777 -4213 5879 -4111
rect 6597 -4213 6699 -4111
<< psubdiff >>
rect -1104 -544 -360 -510
rect -1104 -578 -1070 -544
rect -1036 -578 -1002 -544
rect -968 -578 -934 -544
rect -900 -578 -866 -544
rect -832 -578 -632 -544
rect -598 -578 -564 -544
rect -530 -578 -496 -544
rect -462 -578 -428 -544
rect -394 -578 -360 -544
rect -1104 -611 -360 -578
rect -1104 -612 -1003 -611
rect -1104 -646 -1070 -612
rect -1036 -646 -1003 -612
rect -1104 -680 -1003 -646
rect -461 -612 -360 -611
rect -461 -646 -428 -612
rect -394 -646 -360 -612
rect -1104 -714 -1070 -680
rect -1036 -714 -1003 -680
rect -1104 -748 -1003 -714
rect -1104 -782 -1070 -748
rect -1036 -782 -1003 -748
rect -1104 -982 -1003 -782
rect -1104 -1016 -1070 -982
rect -1036 -1016 -1003 -982
rect -1104 -1050 -1003 -1016
rect -1104 -1084 -1070 -1050
rect -1036 -1084 -1003 -1050
rect -1104 -1118 -1003 -1084
rect -461 -680 -360 -646
rect -461 -714 -428 -680
rect -394 -714 -360 -680
rect -461 -748 -360 -714
rect -461 -782 -428 -748
rect -394 -782 -360 -748
rect -461 -982 -360 -782
rect -461 -1016 -428 -982
rect -394 -1016 -360 -982
rect -461 -1050 -360 -1016
rect -461 -1084 -428 -1050
rect -394 -1084 -360 -1050
rect -1104 -1152 -1070 -1118
rect -1036 -1152 -1003 -1118
rect -1104 -1153 -1003 -1152
rect -461 -1118 -360 -1084
rect -461 -1152 -428 -1118
rect -394 -1152 -360 -1118
rect -461 -1153 -360 -1152
rect -1104 -1186 -360 -1153
rect -1104 -1220 -1070 -1186
rect -1036 -1220 -1002 -1186
rect -968 -1220 -934 -1186
rect -900 -1220 -866 -1186
rect -832 -1220 -632 -1186
rect -598 -1220 -564 -1186
rect -530 -1220 -496 -1186
rect -462 -1220 -428 -1186
rect -394 -1220 -360 -1186
rect -1104 -1254 -360 -1220
rect -284 -544 460 -510
rect -284 -578 -250 -544
rect -216 -578 -182 -544
rect -148 -578 -114 -544
rect -80 -578 -46 -544
rect -12 -578 188 -544
rect 222 -578 256 -544
rect 290 -578 324 -544
rect 358 -578 392 -544
rect 426 -578 460 -544
rect -284 -611 460 -578
rect -284 -612 -183 -611
rect -284 -646 -250 -612
rect -216 -646 -183 -612
rect -284 -680 -183 -646
rect 359 -612 460 -611
rect 359 -646 392 -612
rect 426 -646 460 -612
rect -284 -714 -250 -680
rect -216 -714 -183 -680
rect -284 -748 -183 -714
rect -284 -782 -250 -748
rect -216 -782 -183 -748
rect -284 -982 -183 -782
rect -284 -1016 -250 -982
rect -216 -1016 -183 -982
rect -284 -1050 -183 -1016
rect -284 -1084 -250 -1050
rect -216 -1084 -183 -1050
rect -284 -1118 -183 -1084
rect 359 -680 460 -646
rect 359 -714 392 -680
rect 426 -714 460 -680
rect 359 -748 460 -714
rect 359 -782 392 -748
rect 426 -782 460 -748
rect 359 -982 460 -782
rect 359 -1016 392 -982
rect 426 -1016 460 -982
rect 359 -1050 460 -1016
rect 359 -1084 392 -1050
rect 426 -1084 460 -1050
rect -284 -1152 -250 -1118
rect -216 -1152 -183 -1118
rect -284 -1153 -183 -1152
rect 359 -1118 460 -1084
rect 359 -1152 392 -1118
rect 426 -1152 460 -1118
rect 359 -1153 460 -1152
rect -284 -1186 460 -1153
rect -284 -1220 -250 -1186
rect -216 -1220 -182 -1186
rect -148 -1220 -114 -1186
rect -80 -1220 -46 -1186
rect -12 -1220 188 -1186
rect 222 -1220 256 -1186
rect 290 -1220 324 -1186
rect 358 -1220 392 -1186
rect 426 -1220 460 -1186
rect -284 -1254 460 -1220
rect 536 -544 1280 -510
rect 536 -578 570 -544
rect 604 -578 638 -544
rect 672 -578 706 -544
rect 740 -578 774 -544
rect 808 -578 1008 -544
rect 1042 -578 1076 -544
rect 1110 -578 1144 -544
rect 1178 -578 1212 -544
rect 1246 -578 1280 -544
rect 536 -611 1280 -578
rect 536 -612 637 -611
rect 536 -646 570 -612
rect 604 -646 637 -612
rect 536 -680 637 -646
rect 1179 -612 1280 -611
rect 1179 -646 1212 -612
rect 1246 -646 1280 -612
rect 536 -714 570 -680
rect 604 -714 637 -680
rect 536 -748 637 -714
rect 536 -782 570 -748
rect 604 -782 637 -748
rect 536 -982 637 -782
rect 536 -1016 570 -982
rect 604 -1016 637 -982
rect 536 -1050 637 -1016
rect 536 -1084 570 -1050
rect 604 -1084 637 -1050
rect 536 -1118 637 -1084
rect 1179 -680 1280 -646
rect 1179 -714 1212 -680
rect 1246 -714 1280 -680
rect 1179 -748 1280 -714
rect 1179 -782 1212 -748
rect 1246 -782 1280 -748
rect 1179 -982 1280 -782
rect 1179 -1016 1212 -982
rect 1246 -1016 1280 -982
rect 1179 -1050 1280 -1016
rect 1179 -1084 1212 -1050
rect 1246 -1084 1280 -1050
rect 536 -1152 570 -1118
rect 604 -1152 637 -1118
rect 536 -1153 637 -1152
rect 1179 -1118 1280 -1084
rect 1179 -1152 1212 -1118
rect 1246 -1152 1280 -1118
rect 1179 -1153 1280 -1152
rect 536 -1186 1280 -1153
rect 536 -1220 570 -1186
rect 604 -1220 638 -1186
rect 672 -1220 706 -1186
rect 740 -1220 774 -1186
rect 808 -1220 1008 -1186
rect 1042 -1220 1076 -1186
rect 1110 -1220 1144 -1186
rect 1178 -1220 1212 -1186
rect 1246 -1220 1280 -1186
rect 536 -1254 1280 -1220
rect 1356 -544 2100 -510
rect 1356 -578 1390 -544
rect 1424 -578 1458 -544
rect 1492 -578 1526 -544
rect 1560 -578 1594 -544
rect 1628 -578 1828 -544
rect 1862 -578 1896 -544
rect 1930 -578 1964 -544
rect 1998 -578 2032 -544
rect 2066 -578 2100 -544
rect 1356 -611 2100 -578
rect 1356 -612 1457 -611
rect 1356 -646 1390 -612
rect 1424 -646 1457 -612
rect 1356 -680 1457 -646
rect 1999 -612 2100 -611
rect 1999 -646 2032 -612
rect 2066 -646 2100 -612
rect 1356 -714 1390 -680
rect 1424 -714 1457 -680
rect 1356 -748 1457 -714
rect 1356 -782 1390 -748
rect 1424 -782 1457 -748
rect 1356 -982 1457 -782
rect 1356 -1016 1390 -982
rect 1424 -1016 1457 -982
rect 1356 -1050 1457 -1016
rect 1356 -1084 1390 -1050
rect 1424 -1084 1457 -1050
rect 1356 -1118 1457 -1084
rect 1999 -680 2100 -646
rect 1999 -714 2032 -680
rect 2066 -714 2100 -680
rect 1999 -748 2100 -714
rect 1999 -782 2032 -748
rect 2066 -782 2100 -748
rect 1999 -982 2100 -782
rect 1999 -1016 2032 -982
rect 2066 -1016 2100 -982
rect 1999 -1050 2100 -1016
rect 1999 -1084 2032 -1050
rect 2066 -1084 2100 -1050
rect 1356 -1152 1390 -1118
rect 1424 -1152 1457 -1118
rect 1356 -1153 1457 -1152
rect 1999 -1118 2100 -1084
rect 1999 -1152 2032 -1118
rect 2066 -1152 2100 -1118
rect 1999 -1153 2100 -1152
rect 1356 -1186 2100 -1153
rect 1356 -1220 1390 -1186
rect 1424 -1220 1458 -1186
rect 1492 -1220 1526 -1186
rect 1560 -1220 1594 -1186
rect 1628 -1220 1828 -1186
rect 1862 -1220 1896 -1186
rect 1930 -1220 1964 -1186
rect 1998 -1220 2032 -1186
rect 2066 -1220 2100 -1186
rect 1356 -1254 2100 -1220
rect 2176 -544 2920 -510
rect 2176 -578 2210 -544
rect 2244 -578 2278 -544
rect 2312 -578 2346 -544
rect 2380 -578 2414 -544
rect 2448 -578 2648 -544
rect 2682 -578 2716 -544
rect 2750 -578 2784 -544
rect 2818 -578 2852 -544
rect 2886 -578 2920 -544
rect 2176 -611 2920 -578
rect 2176 -612 2277 -611
rect 2176 -646 2210 -612
rect 2244 -646 2277 -612
rect 2176 -680 2277 -646
rect 2819 -612 2920 -611
rect 2819 -646 2852 -612
rect 2886 -646 2920 -612
rect 2176 -714 2210 -680
rect 2244 -714 2277 -680
rect 2176 -748 2277 -714
rect 2176 -782 2210 -748
rect 2244 -782 2277 -748
rect 2176 -982 2277 -782
rect 2176 -1016 2210 -982
rect 2244 -1016 2277 -982
rect 2176 -1050 2277 -1016
rect 2176 -1084 2210 -1050
rect 2244 -1084 2277 -1050
rect 2176 -1118 2277 -1084
rect 2819 -680 2920 -646
rect 2819 -714 2852 -680
rect 2886 -714 2920 -680
rect 2819 -748 2920 -714
rect 2819 -782 2852 -748
rect 2886 -782 2920 -748
rect 2819 -982 2920 -782
rect 2819 -1016 2852 -982
rect 2886 -1016 2920 -982
rect 2819 -1050 2920 -1016
rect 2819 -1084 2852 -1050
rect 2886 -1084 2920 -1050
rect 2176 -1152 2210 -1118
rect 2244 -1152 2277 -1118
rect 2176 -1153 2277 -1152
rect 2819 -1118 2920 -1084
rect 2819 -1152 2852 -1118
rect 2886 -1152 2920 -1118
rect 2819 -1153 2920 -1152
rect 2176 -1186 2920 -1153
rect 2176 -1220 2210 -1186
rect 2244 -1220 2278 -1186
rect 2312 -1220 2346 -1186
rect 2380 -1220 2414 -1186
rect 2448 -1220 2648 -1186
rect 2682 -1220 2716 -1186
rect 2750 -1220 2784 -1186
rect 2818 -1220 2852 -1186
rect 2886 -1220 2920 -1186
rect 2176 -1254 2920 -1220
rect 2996 -544 3740 -510
rect 2996 -578 3030 -544
rect 3064 -578 3098 -544
rect 3132 -578 3166 -544
rect 3200 -578 3234 -544
rect 3268 -578 3468 -544
rect 3502 -578 3536 -544
rect 3570 -578 3604 -544
rect 3638 -578 3672 -544
rect 3706 -578 3740 -544
rect 2996 -611 3740 -578
rect 2996 -612 3097 -611
rect 2996 -646 3030 -612
rect 3064 -646 3097 -612
rect 2996 -680 3097 -646
rect 3639 -612 3740 -611
rect 3639 -646 3672 -612
rect 3706 -646 3740 -612
rect 2996 -714 3030 -680
rect 3064 -714 3097 -680
rect 2996 -748 3097 -714
rect 2996 -782 3030 -748
rect 3064 -782 3097 -748
rect 2996 -982 3097 -782
rect 2996 -1016 3030 -982
rect 3064 -1016 3097 -982
rect 2996 -1050 3097 -1016
rect 2996 -1084 3030 -1050
rect 3064 -1084 3097 -1050
rect 2996 -1118 3097 -1084
rect 3639 -680 3740 -646
rect 3639 -714 3672 -680
rect 3706 -714 3740 -680
rect 3639 -748 3740 -714
rect 3639 -782 3672 -748
rect 3706 -782 3740 -748
rect 3639 -982 3740 -782
rect 3639 -1016 3672 -982
rect 3706 -1016 3740 -982
rect 3639 -1050 3740 -1016
rect 3639 -1084 3672 -1050
rect 3706 -1084 3740 -1050
rect 2996 -1152 3030 -1118
rect 3064 -1152 3097 -1118
rect 2996 -1153 3097 -1152
rect 3639 -1118 3740 -1084
rect 3639 -1152 3672 -1118
rect 3706 -1152 3740 -1118
rect 3639 -1153 3740 -1152
rect 2996 -1186 3740 -1153
rect 2996 -1220 3030 -1186
rect 3064 -1220 3098 -1186
rect 3132 -1220 3166 -1186
rect 3200 -1220 3234 -1186
rect 3268 -1220 3468 -1186
rect 3502 -1220 3536 -1186
rect 3570 -1220 3604 -1186
rect 3638 -1220 3672 -1186
rect 3706 -1220 3740 -1186
rect 2996 -1254 3740 -1220
rect 3816 -544 4560 -510
rect 3816 -578 3850 -544
rect 3884 -578 3918 -544
rect 3952 -578 3986 -544
rect 4020 -578 4054 -544
rect 4088 -578 4288 -544
rect 4322 -578 4356 -544
rect 4390 -578 4424 -544
rect 4458 -578 4492 -544
rect 4526 -578 4560 -544
rect 3816 -611 4560 -578
rect 3816 -612 3917 -611
rect 3816 -646 3850 -612
rect 3884 -646 3917 -612
rect 3816 -680 3917 -646
rect 4459 -612 4560 -611
rect 4459 -646 4492 -612
rect 4526 -646 4560 -612
rect 3816 -714 3850 -680
rect 3884 -714 3917 -680
rect 3816 -748 3917 -714
rect 3816 -782 3850 -748
rect 3884 -782 3917 -748
rect 3816 -982 3917 -782
rect 3816 -1016 3850 -982
rect 3884 -1016 3917 -982
rect 3816 -1050 3917 -1016
rect 3816 -1084 3850 -1050
rect 3884 -1084 3917 -1050
rect 3816 -1118 3917 -1084
rect 4459 -680 4560 -646
rect 4459 -714 4492 -680
rect 4526 -714 4560 -680
rect 4459 -748 4560 -714
rect 4459 -782 4492 -748
rect 4526 -782 4560 -748
rect 4459 -982 4560 -782
rect 4459 -1016 4492 -982
rect 4526 -1016 4560 -982
rect 4459 -1050 4560 -1016
rect 4459 -1084 4492 -1050
rect 4526 -1084 4560 -1050
rect 3816 -1152 3850 -1118
rect 3884 -1152 3917 -1118
rect 3816 -1153 3917 -1152
rect 4459 -1118 4560 -1084
rect 4459 -1152 4492 -1118
rect 4526 -1152 4560 -1118
rect 4459 -1153 4560 -1152
rect 3816 -1186 4560 -1153
rect 3816 -1220 3850 -1186
rect 3884 -1220 3918 -1186
rect 3952 -1220 3986 -1186
rect 4020 -1220 4054 -1186
rect 4088 -1220 4288 -1186
rect 4322 -1220 4356 -1186
rect 4390 -1220 4424 -1186
rect 4458 -1220 4492 -1186
rect 4526 -1220 4560 -1186
rect 3816 -1254 4560 -1220
rect 4636 -544 5380 -510
rect 4636 -578 4670 -544
rect 4704 -578 4738 -544
rect 4772 -578 4806 -544
rect 4840 -578 4874 -544
rect 4908 -578 5108 -544
rect 5142 -578 5176 -544
rect 5210 -578 5244 -544
rect 5278 -578 5312 -544
rect 5346 -578 5380 -544
rect 4636 -611 5380 -578
rect 4636 -612 4737 -611
rect 4636 -646 4670 -612
rect 4704 -646 4737 -612
rect 4636 -680 4737 -646
rect 5279 -612 5380 -611
rect 5279 -646 5312 -612
rect 5346 -646 5380 -612
rect 4636 -714 4670 -680
rect 4704 -714 4737 -680
rect 4636 -748 4737 -714
rect 4636 -782 4670 -748
rect 4704 -782 4737 -748
rect 4636 -982 4737 -782
rect 4636 -1016 4670 -982
rect 4704 -1016 4737 -982
rect 4636 -1050 4737 -1016
rect 4636 -1084 4670 -1050
rect 4704 -1084 4737 -1050
rect 4636 -1118 4737 -1084
rect 5279 -680 5380 -646
rect 5279 -714 5312 -680
rect 5346 -714 5380 -680
rect 5279 -748 5380 -714
rect 5279 -782 5312 -748
rect 5346 -782 5380 -748
rect 5279 -982 5380 -782
rect 5279 -1016 5312 -982
rect 5346 -1016 5380 -982
rect 5279 -1050 5380 -1016
rect 5279 -1084 5312 -1050
rect 5346 -1084 5380 -1050
rect 4636 -1152 4670 -1118
rect 4704 -1152 4737 -1118
rect 4636 -1153 4737 -1152
rect 5279 -1118 5380 -1084
rect 5279 -1152 5312 -1118
rect 5346 -1152 5380 -1118
rect 5279 -1153 5380 -1152
rect 4636 -1186 5380 -1153
rect 4636 -1220 4670 -1186
rect 4704 -1220 4738 -1186
rect 4772 -1220 4806 -1186
rect 4840 -1220 4874 -1186
rect 4908 -1220 5108 -1186
rect 5142 -1220 5176 -1186
rect 5210 -1220 5244 -1186
rect 5278 -1220 5312 -1186
rect 5346 -1220 5380 -1186
rect 4636 -1254 5380 -1220
rect 5456 -544 6200 -510
rect 5456 -578 5490 -544
rect 5524 -578 5558 -544
rect 5592 -578 5626 -544
rect 5660 -578 5694 -544
rect 5728 -578 5928 -544
rect 5962 -578 5996 -544
rect 6030 -578 6064 -544
rect 6098 -578 6132 -544
rect 6166 -578 6200 -544
rect 5456 -611 6200 -578
rect 5456 -612 5557 -611
rect 5456 -646 5490 -612
rect 5524 -646 5557 -612
rect 5456 -680 5557 -646
rect 6099 -612 6200 -611
rect 6099 -646 6132 -612
rect 6166 -646 6200 -612
rect 5456 -714 5490 -680
rect 5524 -714 5557 -680
rect 5456 -748 5557 -714
rect 5456 -782 5490 -748
rect 5524 -782 5557 -748
rect 5456 -982 5557 -782
rect 5456 -1016 5490 -982
rect 5524 -1016 5557 -982
rect 5456 -1050 5557 -1016
rect 5456 -1084 5490 -1050
rect 5524 -1084 5557 -1050
rect 5456 -1118 5557 -1084
rect 6099 -680 6200 -646
rect 6099 -714 6132 -680
rect 6166 -714 6200 -680
rect 6099 -748 6200 -714
rect 6099 -782 6132 -748
rect 6166 -782 6200 -748
rect 6099 -982 6200 -782
rect 6099 -1016 6132 -982
rect 6166 -1016 6200 -982
rect 6099 -1050 6200 -1016
rect 6099 -1084 6132 -1050
rect 6166 -1084 6200 -1050
rect 5456 -1152 5490 -1118
rect 5524 -1152 5557 -1118
rect 5456 -1153 5557 -1152
rect 6099 -1118 6200 -1084
rect 6099 -1152 6132 -1118
rect 6166 -1152 6200 -1118
rect 6099 -1153 6200 -1152
rect 5456 -1186 6200 -1153
rect 5456 -1220 5490 -1186
rect 5524 -1220 5558 -1186
rect 5592 -1220 5626 -1186
rect 5660 -1220 5694 -1186
rect 5728 -1220 5928 -1186
rect 5962 -1220 5996 -1186
rect 6030 -1220 6064 -1186
rect 6098 -1220 6132 -1186
rect 6166 -1220 6200 -1186
rect 5456 -1254 6200 -1220
rect 6276 -544 7020 -510
rect 6276 -578 6310 -544
rect 6344 -578 6378 -544
rect 6412 -578 6446 -544
rect 6480 -578 6514 -544
rect 6548 -578 6748 -544
rect 6782 -578 6816 -544
rect 6850 -578 6884 -544
rect 6918 -578 6952 -544
rect 6986 -578 7020 -544
rect 6276 -611 7020 -578
rect 6276 -612 6377 -611
rect 6276 -646 6310 -612
rect 6344 -646 6377 -612
rect 6276 -680 6377 -646
rect 6919 -612 7020 -611
rect 6919 -646 6952 -612
rect 6986 -646 7020 -612
rect 6276 -714 6310 -680
rect 6344 -714 6377 -680
rect 6276 -748 6377 -714
rect 6276 -782 6310 -748
rect 6344 -782 6377 -748
rect 6276 -982 6377 -782
rect 6276 -1016 6310 -982
rect 6344 -1016 6377 -982
rect 6276 -1050 6377 -1016
rect 6276 -1084 6310 -1050
rect 6344 -1084 6377 -1050
rect 6276 -1118 6377 -1084
rect 6919 -680 7020 -646
rect 6919 -714 6952 -680
rect 6986 -714 7020 -680
rect 6919 -748 7020 -714
rect 6919 -782 6952 -748
rect 6986 -782 7020 -748
rect 6919 -982 7020 -782
rect 6919 -1016 6952 -982
rect 6986 -1016 7020 -982
rect 6919 -1050 7020 -1016
rect 6919 -1084 6952 -1050
rect 6986 -1084 7020 -1050
rect 6276 -1152 6310 -1118
rect 6344 -1152 6377 -1118
rect 6276 -1153 6377 -1152
rect 6919 -1118 7020 -1084
rect 6919 -1152 6952 -1118
rect 6986 -1152 7020 -1118
rect 6919 -1153 7020 -1152
rect 6276 -1186 7020 -1153
rect 6276 -1220 6310 -1186
rect 6344 -1220 6378 -1186
rect 6412 -1220 6446 -1186
rect 6480 -1220 6514 -1186
rect 6548 -1220 6748 -1186
rect 6782 -1220 6816 -1186
rect 6850 -1220 6884 -1186
rect 6918 -1220 6952 -1186
rect 6986 -1220 7020 -1186
rect 6276 -1254 7020 -1220
rect 7126 -544 7870 -510
rect 7126 -578 7160 -544
rect 7194 -578 7228 -544
rect 7262 -578 7296 -544
rect 7330 -578 7364 -544
rect 7398 -578 7598 -544
rect 7632 -578 7666 -544
rect 7700 -578 7734 -544
rect 7768 -578 7802 -544
rect 7836 -578 7870 -544
rect 7126 -611 7870 -578
rect 7126 -612 7227 -611
rect 7126 -646 7160 -612
rect 7194 -646 7227 -612
rect 7126 -680 7227 -646
rect 7769 -612 7870 -611
rect 7769 -646 7802 -612
rect 7836 -646 7870 -612
rect 7126 -714 7160 -680
rect 7194 -714 7227 -680
rect 7126 -748 7227 -714
rect 7126 -782 7160 -748
rect 7194 -782 7227 -748
rect 7126 -982 7227 -782
rect 7126 -1016 7160 -982
rect 7194 -1016 7227 -982
rect 7126 -1050 7227 -1016
rect 7126 -1084 7160 -1050
rect 7194 -1084 7227 -1050
rect 7126 -1118 7227 -1084
rect 7769 -680 7870 -646
rect 7769 -714 7802 -680
rect 7836 -714 7870 -680
rect 7769 -748 7870 -714
rect 7769 -782 7802 -748
rect 7836 -782 7870 -748
rect 7769 -982 7870 -782
rect 7769 -1016 7802 -982
rect 7836 -1016 7870 -982
rect 7769 -1050 7870 -1016
rect 7769 -1084 7802 -1050
rect 7836 -1084 7870 -1050
rect 7126 -1152 7160 -1118
rect 7194 -1152 7227 -1118
rect 7126 -1153 7227 -1152
rect 7769 -1118 7870 -1084
rect 7769 -1152 7802 -1118
rect 7836 -1152 7870 -1118
rect 7769 -1153 7870 -1152
rect 7126 -1186 7870 -1153
rect 7126 -1220 7160 -1186
rect 7194 -1220 7228 -1186
rect 7262 -1220 7296 -1186
rect 7330 -1220 7364 -1186
rect 7398 -1220 7598 -1186
rect 7632 -1220 7666 -1186
rect 7700 -1220 7734 -1186
rect 7768 -1220 7802 -1186
rect 7836 -1220 7870 -1186
rect 7126 -1254 7870 -1220
rect -1104 -1364 -360 -1330
rect -1104 -1398 -1070 -1364
rect -1036 -1398 -1002 -1364
rect -968 -1398 -934 -1364
rect -900 -1398 -866 -1364
rect -832 -1398 -632 -1364
rect -598 -1398 -564 -1364
rect -530 -1398 -496 -1364
rect -462 -1398 -428 -1364
rect -394 -1398 -360 -1364
rect -1104 -1431 -360 -1398
rect -1104 -1432 -1003 -1431
rect -1104 -1466 -1070 -1432
rect -1036 -1466 -1003 -1432
rect -1104 -1500 -1003 -1466
rect -461 -1432 -360 -1431
rect -461 -1466 -428 -1432
rect -394 -1466 -360 -1432
rect -1104 -1534 -1070 -1500
rect -1036 -1534 -1003 -1500
rect -1104 -1568 -1003 -1534
rect -1104 -1602 -1070 -1568
rect -1036 -1602 -1003 -1568
rect -1104 -1802 -1003 -1602
rect -1104 -1836 -1070 -1802
rect -1036 -1836 -1003 -1802
rect -1104 -1870 -1003 -1836
rect -1104 -1904 -1070 -1870
rect -1036 -1904 -1003 -1870
rect -1104 -1938 -1003 -1904
rect -461 -1500 -360 -1466
rect -461 -1534 -428 -1500
rect -394 -1534 -360 -1500
rect -461 -1568 -360 -1534
rect -461 -1602 -428 -1568
rect -394 -1602 -360 -1568
rect -461 -1802 -360 -1602
rect -461 -1836 -428 -1802
rect -394 -1836 -360 -1802
rect -461 -1870 -360 -1836
rect -461 -1904 -428 -1870
rect -394 -1904 -360 -1870
rect -1104 -1972 -1070 -1938
rect -1036 -1972 -1003 -1938
rect -1104 -1973 -1003 -1972
rect -461 -1938 -360 -1904
rect -461 -1972 -428 -1938
rect -394 -1972 -360 -1938
rect -461 -1973 -360 -1972
rect -1104 -2006 -360 -1973
rect -1104 -2040 -1070 -2006
rect -1036 -2040 -1002 -2006
rect -968 -2040 -934 -2006
rect -900 -2040 -866 -2006
rect -832 -2040 -632 -2006
rect -598 -2040 -564 -2006
rect -530 -2040 -496 -2006
rect -462 -2040 -428 -2006
rect -394 -2040 -360 -2006
rect -1104 -2074 -360 -2040
rect -284 -1364 460 -1330
rect -284 -1398 -250 -1364
rect -216 -1398 -182 -1364
rect -148 -1398 -114 -1364
rect -80 -1398 -46 -1364
rect -12 -1398 188 -1364
rect 222 -1398 256 -1364
rect 290 -1398 324 -1364
rect 358 -1398 392 -1364
rect 426 -1398 460 -1364
rect -284 -1431 460 -1398
rect -284 -1432 -183 -1431
rect -284 -1466 -250 -1432
rect -216 -1466 -183 -1432
rect -284 -1500 -183 -1466
rect 359 -1432 460 -1431
rect 359 -1466 392 -1432
rect 426 -1466 460 -1432
rect -284 -1534 -250 -1500
rect -216 -1534 -183 -1500
rect -284 -1568 -183 -1534
rect -284 -1602 -250 -1568
rect -216 -1602 -183 -1568
rect -284 -1802 -183 -1602
rect -284 -1836 -250 -1802
rect -216 -1836 -183 -1802
rect -284 -1870 -183 -1836
rect -284 -1904 -250 -1870
rect -216 -1904 -183 -1870
rect -284 -1938 -183 -1904
rect 359 -1500 460 -1466
rect 359 -1534 392 -1500
rect 426 -1534 460 -1500
rect 359 -1568 460 -1534
rect 359 -1602 392 -1568
rect 426 -1602 460 -1568
rect 359 -1802 460 -1602
rect 359 -1836 392 -1802
rect 426 -1836 460 -1802
rect 359 -1870 460 -1836
rect 359 -1904 392 -1870
rect 426 -1904 460 -1870
rect -284 -1972 -250 -1938
rect -216 -1972 -183 -1938
rect -284 -1973 -183 -1972
rect 359 -1938 460 -1904
rect 359 -1972 392 -1938
rect 426 -1972 460 -1938
rect 359 -1973 460 -1972
rect -284 -2006 460 -1973
rect -284 -2040 -250 -2006
rect -216 -2040 -182 -2006
rect -148 -2040 -114 -2006
rect -80 -2040 -46 -2006
rect -12 -2040 188 -2006
rect 222 -2040 256 -2006
rect 290 -2040 324 -2006
rect 358 -2040 392 -2006
rect 426 -2040 460 -2006
rect -284 -2074 460 -2040
rect 536 -1364 1280 -1330
rect 536 -1398 570 -1364
rect 604 -1398 638 -1364
rect 672 -1398 706 -1364
rect 740 -1398 774 -1364
rect 808 -1398 1008 -1364
rect 1042 -1398 1076 -1364
rect 1110 -1398 1144 -1364
rect 1178 -1398 1212 -1364
rect 1246 -1398 1280 -1364
rect 536 -1431 1280 -1398
rect 536 -1432 637 -1431
rect 536 -1466 570 -1432
rect 604 -1466 637 -1432
rect 536 -1500 637 -1466
rect 1179 -1432 1280 -1431
rect 1179 -1466 1212 -1432
rect 1246 -1466 1280 -1432
rect 536 -1534 570 -1500
rect 604 -1534 637 -1500
rect 536 -1568 637 -1534
rect 536 -1602 570 -1568
rect 604 -1602 637 -1568
rect 536 -1802 637 -1602
rect 536 -1836 570 -1802
rect 604 -1836 637 -1802
rect 536 -1870 637 -1836
rect 536 -1904 570 -1870
rect 604 -1904 637 -1870
rect 536 -1938 637 -1904
rect 1179 -1500 1280 -1466
rect 1179 -1534 1212 -1500
rect 1246 -1534 1280 -1500
rect 1179 -1568 1280 -1534
rect 1179 -1602 1212 -1568
rect 1246 -1602 1280 -1568
rect 1179 -1802 1280 -1602
rect 1179 -1836 1212 -1802
rect 1246 -1836 1280 -1802
rect 1179 -1870 1280 -1836
rect 1179 -1904 1212 -1870
rect 1246 -1904 1280 -1870
rect 536 -1972 570 -1938
rect 604 -1972 637 -1938
rect 536 -1973 637 -1972
rect 1179 -1938 1280 -1904
rect 1179 -1972 1212 -1938
rect 1246 -1972 1280 -1938
rect 1179 -1973 1280 -1972
rect 536 -2006 1280 -1973
rect 536 -2040 570 -2006
rect 604 -2040 638 -2006
rect 672 -2040 706 -2006
rect 740 -2040 774 -2006
rect 808 -2040 1008 -2006
rect 1042 -2040 1076 -2006
rect 1110 -2040 1144 -2006
rect 1178 -2040 1212 -2006
rect 1246 -2040 1280 -2006
rect 536 -2074 1280 -2040
rect 1356 -1364 2100 -1330
rect 1356 -1398 1390 -1364
rect 1424 -1398 1458 -1364
rect 1492 -1398 1526 -1364
rect 1560 -1398 1594 -1364
rect 1628 -1398 1828 -1364
rect 1862 -1398 1896 -1364
rect 1930 -1398 1964 -1364
rect 1998 -1398 2032 -1364
rect 2066 -1398 2100 -1364
rect 1356 -1431 2100 -1398
rect 1356 -1432 1457 -1431
rect 1356 -1466 1390 -1432
rect 1424 -1466 1457 -1432
rect 1356 -1500 1457 -1466
rect 1999 -1432 2100 -1431
rect 1999 -1466 2032 -1432
rect 2066 -1466 2100 -1432
rect 1356 -1534 1390 -1500
rect 1424 -1534 1457 -1500
rect 1356 -1568 1457 -1534
rect 1356 -1602 1390 -1568
rect 1424 -1602 1457 -1568
rect 1356 -1802 1457 -1602
rect 1356 -1836 1390 -1802
rect 1424 -1836 1457 -1802
rect 1356 -1870 1457 -1836
rect 1356 -1904 1390 -1870
rect 1424 -1904 1457 -1870
rect 1356 -1938 1457 -1904
rect 1999 -1500 2100 -1466
rect 1999 -1534 2032 -1500
rect 2066 -1534 2100 -1500
rect 1999 -1568 2100 -1534
rect 1999 -1602 2032 -1568
rect 2066 -1602 2100 -1568
rect 1999 -1802 2100 -1602
rect 1999 -1836 2032 -1802
rect 2066 -1836 2100 -1802
rect 1999 -1870 2100 -1836
rect 1999 -1904 2032 -1870
rect 2066 -1904 2100 -1870
rect 1356 -1972 1390 -1938
rect 1424 -1972 1457 -1938
rect 1356 -1973 1457 -1972
rect 1999 -1938 2100 -1904
rect 1999 -1972 2032 -1938
rect 2066 -1972 2100 -1938
rect 1999 -1973 2100 -1972
rect 1356 -2006 2100 -1973
rect 1356 -2040 1390 -2006
rect 1424 -2040 1458 -2006
rect 1492 -2040 1526 -2006
rect 1560 -2040 1594 -2006
rect 1628 -2040 1828 -2006
rect 1862 -2040 1896 -2006
rect 1930 -2040 1964 -2006
rect 1998 -2040 2032 -2006
rect 2066 -2040 2100 -2006
rect 1356 -2074 2100 -2040
rect 2176 -1364 2920 -1330
rect 2176 -1398 2210 -1364
rect 2244 -1398 2278 -1364
rect 2312 -1398 2346 -1364
rect 2380 -1398 2414 -1364
rect 2448 -1398 2648 -1364
rect 2682 -1398 2716 -1364
rect 2750 -1398 2784 -1364
rect 2818 -1398 2852 -1364
rect 2886 -1398 2920 -1364
rect 2176 -1431 2920 -1398
rect 2176 -1432 2277 -1431
rect 2176 -1466 2210 -1432
rect 2244 -1466 2277 -1432
rect 2176 -1500 2277 -1466
rect 2819 -1432 2920 -1431
rect 2819 -1466 2852 -1432
rect 2886 -1466 2920 -1432
rect 2176 -1534 2210 -1500
rect 2244 -1534 2277 -1500
rect 2176 -1568 2277 -1534
rect 2176 -1602 2210 -1568
rect 2244 -1602 2277 -1568
rect 2176 -1802 2277 -1602
rect 2176 -1836 2210 -1802
rect 2244 -1836 2277 -1802
rect 2176 -1870 2277 -1836
rect 2176 -1904 2210 -1870
rect 2244 -1904 2277 -1870
rect 2176 -1938 2277 -1904
rect 2819 -1500 2920 -1466
rect 2819 -1534 2852 -1500
rect 2886 -1534 2920 -1500
rect 2819 -1568 2920 -1534
rect 2819 -1602 2852 -1568
rect 2886 -1602 2920 -1568
rect 2819 -1802 2920 -1602
rect 2819 -1836 2852 -1802
rect 2886 -1836 2920 -1802
rect 2819 -1870 2920 -1836
rect 2819 -1904 2852 -1870
rect 2886 -1904 2920 -1870
rect 2176 -1972 2210 -1938
rect 2244 -1972 2277 -1938
rect 2176 -1973 2277 -1972
rect 2819 -1938 2920 -1904
rect 2819 -1972 2852 -1938
rect 2886 -1972 2920 -1938
rect 2819 -1973 2920 -1972
rect 2176 -2006 2920 -1973
rect 2176 -2040 2210 -2006
rect 2244 -2040 2278 -2006
rect 2312 -2040 2346 -2006
rect 2380 -2040 2414 -2006
rect 2448 -2040 2648 -2006
rect 2682 -2040 2716 -2006
rect 2750 -2040 2784 -2006
rect 2818 -2040 2852 -2006
rect 2886 -2040 2920 -2006
rect 2176 -2074 2920 -2040
rect 2996 -1364 3740 -1330
rect 2996 -1398 3030 -1364
rect 3064 -1398 3098 -1364
rect 3132 -1398 3166 -1364
rect 3200 -1398 3234 -1364
rect 3268 -1398 3468 -1364
rect 3502 -1398 3536 -1364
rect 3570 -1398 3604 -1364
rect 3638 -1398 3672 -1364
rect 3706 -1398 3740 -1364
rect 2996 -1431 3740 -1398
rect 2996 -1432 3097 -1431
rect 2996 -1466 3030 -1432
rect 3064 -1466 3097 -1432
rect 2996 -1500 3097 -1466
rect 3639 -1432 3740 -1431
rect 3639 -1466 3672 -1432
rect 3706 -1466 3740 -1432
rect 2996 -1534 3030 -1500
rect 3064 -1534 3097 -1500
rect 2996 -1568 3097 -1534
rect 2996 -1602 3030 -1568
rect 3064 -1602 3097 -1568
rect 2996 -1802 3097 -1602
rect 2996 -1836 3030 -1802
rect 3064 -1836 3097 -1802
rect 2996 -1870 3097 -1836
rect 2996 -1904 3030 -1870
rect 3064 -1904 3097 -1870
rect 2996 -1938 3097 -1904
rect 3639 -1500 3740 -1466
rect 3639 -1534 3672 -1500
rect 3706 -1534 3740 -1500
rect 3639 -1568 3740 -1534
rect 3639 -1602 3672 -1568
rect 3706 -1602 3740 -1568
rect 3639 -1802 3740 -1602
rect 3639 -1836 3672 -1802
rect 3706 -1836 3740 -1802
rect 3639 -1870 3740 -1836
rect 3639 -1904 3672 -1870
rect 3706 -1904 3740 -1870
rect 2996 -1972 3030 -1938
rect 3064 -1972 3097 -1938
rect 2996 -1973 3097 -1972
rect 3639 -1938 3740 -1904
rect 3639 -1972 3672 -1938
rect 3706 -1972 3740 -1938
rect 3639 -1973 3740 -1972
rect 2996 -2006 3740 -1973
rect 2996 -2040 3030 -2006
rect 3064 -2040 3098 -2006
rect 3132 -2040 3166 -2006
rect 3200 -2040 3234 -2006
rect 3268 -2040 3468 -2006
rect 3502 -2040 3536 -2006
rect 3570 -2040 3604 -2006
rect 3638 -2040 3672 -2006
rect 3706 -2040 3740 -2006
rect 2996 -2074 3740 -2040
rect 3816 -1364 4560 -1330
rect 3816 -1398 3850 -1364
rect 3884 -1398 3918 -1364
rect 3952 -1398 3986 -1364
rect 4020 -1398 4054 -1364
rect 4088 -1398 4288 -1364
rect 4322 -1398 4356 -1364
rect 4390 -1398 4424 -1364
rect 4458 -1398 4492 -1364
rect 4526 -1398 4560 -1364
rect 3816 -1431 4560 -1398
rect 3816 -1432 3917 -1431
rect 3816 -1466 3850 -1432
rect 3884 -1466 3917 -1432
rect 3816 -1500 3917 -1466
rect 4459 -1432 4560 -1431
rect 4459 -1466 4492 -1432
rect 4526 -1466 4560 -1432
rect 3816 -1534 3850 -1500
rect 3884 -1534 3917 -1500
rect 3816 -1568 3917 -1534
rect 3816 -1602 3850 -1568
rect 3884 -1602 3917 -1568
rect 3816 -1802 3917 -1602
rect 3816 -1836 3850 -1802
rect 3884 -1836 3917 -1802
rect 3816 -1870 3917 -1836
rect 3816 -1904 3850 -1870
rect 3884 -1904 3917 -1870
rect 3816 -1938 3917 -1904
rect 4459 -1500 4560 -1466
rect 4459 -1534 4492 -1500
rect 4526 -1534 4560 -1500
rect 4459 -1568 4560 -1534
rect 4459 -1602 4492 -1568
rect 4526 -1602 4560 -1568
rect 4459 -1802 4560 -1602
rect 4459 -1836 4492 -1802
rect 4526 -1836 4560 -1802
rect 4459 -1870 4560 -1836
rect 4459 -1904 4492 -1870
rect 4526 -1904 4560 -1870
rect 3816 -1972 3850 -1938
rect 3884 -1972 3917 -1938
rect 3816 -1973 3917 -1972
rect 4459 -1938 4560 -1904
rect 4459 -1972 4492 -1938
rect 4526 -1972 4560 -1938
rect 4459 -1973 4560 -1972
rect 3816 -2006 4560 -1973
rect 3816 -2040 3850 -2006
rect 3884 -2040 3918 -2006
rect 3952 -2040 3986 -2006
rect 4020 -2040 4054 -2006
rect 4088 -2040 4288 -2006
rect 4322 -2040 4356 -2006
rect 4390 -2040 4424 -2006
rect 4458 -2040 4492 -2006
rect 4526 -2040 4560 -2006
rect 3816 -2074 4560 -2040
rect 4636 -1364 5380 -1330
rect 4636 -1398 4670 -1364
rect 4704 -1398 4738 -1364
rect 4772 -1398 4806 -1364
rect 4840 -1398 4874 -1364
rect 4908 -1398 5108 -1364
rect 5142 -1398 5176 -1364
rect 5210 -1398 5244 -1364
rect 5278 -1398 5312 -1364
rect 5346 -1398 5380 -1364
rect 4636 -1431 5380 -1398
rect 4636 -1432 4737 -1431
rect 4636 -1466 4670 -1432
rect 4704 -1466 4737 -1432
rect 4636 -1500 4737 -1466
rect 5279 -1432 5380 -1431
rect 5279 -1466 5312 -1432
rect 5346 -1466 5380 -1432
rect 4636 -1534 4670 -1500
rect 4704 -1534 4737 -1500
rect 4636 -1568 4737 -1534
rect 4636 -1602 4670 -1568
rect 4704 -1602 4737 -1568
rect 4636 -1802 4737 -1602
rect 4636 -1836 4670 -1802
rect 4704 -1836 4737 -1802
rect 4636 -1870 4737 -1836
rect 4636 -1904 4670 -1870
rect 4704 -1904 4737 -1870
rect 4636 -1938 4737 -1904
rect 5279 -1500 5380 -1466
rect 5279 -1534 5312 -1500
rect 5346 -1534 5380 -1500
rect 5279 -1568 5380 -1534
rect 5279 -1602 5312 -1568
rect 5346 -1602 5380 -1568
rect 5279 -1802 5380 -1602
rect 5279 -1836 5312 -1802
rect 5346 -1836 5380 -1802
rect 5279 -1870 5380 -1836
rect 5279 -1904 5312 -1870
rect 5346 -1904 5380 -1870
rect 4636 -1972 4670 -1938
rect 4704 -1972 4737 -1938
rect 4636 -1973 4737 -1972
rect 5279 -1938 5380 -1904
rect 5279 -1972 5312 -1938
rect 5346 -1972 5380 -1938
rect 5279 -1973 5380 -1972
rect 4636 -2006 5380 -1973
rect 4636 -2040 4670 -2006
rect 4704 -2040 4738 -2006
rect 4772 -2040 4806 -2006
rect 4840 -2040 4874 -2006
rect 4908 -2040 5108 -2006
rect 5142 -2040 5176 -2006
rect 5210 -2040 5244 -2006
rect 5278 -2040 5312 -2006
rect 5346 -2040 5380 -2006
rect 4636 -2074 5380 -2040
rect 5456 -1364 6200 -1330
rect 5456 -1398 5490 -1364
rect 5524 -1398 5558 -1364
rect 5592 -1398 5626 -1364
rect 5660 -1398 5694 -1364
rect 5728 -1398 5928 -1364
rect 5962 -1398 5996 -1364
rect 6030 -1398 6064 -1364
rect 6098 -1398 6132 -1364
rect 6166 -1398 6200 -1364
rect 5456 -1431 6200 -1398
rect 5456 -1432 5557 -1431
rect 5456 -1466 5490 -1432
rect 5524 -1466 5557 -1432
rect 5456 -1500 5557 -1466
rect 6099 -1432 6200 -1431
rect 6099 -1466 6132 -1432
rect 6166 -1466 6200 -1432
rect 5456 -1534 5490 -1500
rect 5524 -1534 5557 -1500
rect 5456 -1568 5557 -1534
rect 5456 -1602 5490 -1568
rect 5524 -1602 5557 -1568
rect 5456 -1802 5557 -1602
rect 5456 -1836 5490 -1802
rect 5524 -1836 5557 -1802
rect 5456 -1870 5557 -1836
rect 5456 -1904 5490 -1870
rect 5524 -1904 5557 -1870
rect 5456 -1938 5557 -1904
rect 6099 -1500 6200 -1466
rect 6099 -1534 6132 -1500
rect 6166 -1534 6200 -1500
rect 6099 -1568 6200 -1534
rect 6099 -1602 6132 -1568
rect 6166 -1602 6200 -1568
rect 6099 -1802 6200 -1602
rect 6099 -1836 6132 -1802
rect 6166 -1836 6200 -1802
rect 6099 -1870 6200 -1836
rect 6099 -1904 6132 -1870
rect 6166 -1904 6200 -1870
rect 5456 -1972 5490 -1938
rect 5524 -1972 5557 -1938
rect 5456 -1973 5557 -1972
rect 6099 -1938 6200 -1904
rect 6099 -1972 6132 -1938
rect 6166 -1972 6200 -1938
rect 6099 -1973 6200 -1972
rect 5456 -2006 6200 -1973
rect 5456 -2040 5490 -2006
rect 5524 -2040 5558 -2006
rect 5592 -2040 5626 -2006
rect 5660 -2040 5694 -2006
rect 5728 -2040 5928 -2006
rect 5962 -2040 5996 -2006
rect 6030 -2040 6064 -2006
rect 6098 -2040 6132 -2006
rect 6166 -2040 6200 -2006
rect 5456 -2074 6200 -2040
rect 6276 -1364 7020 -1330
rect 6276 -1398 6310 -1364
rect 6344 -1398 6378 -1364
rect 6412 -1398 6446 -1364
rect 6480 -1398 6514 -1364
rect 6548 -1398 6748 -1364
rect 6782 -1398 6816 -1364
rect 6850 -1398 6884 -1364
rect 6918 -1398 6952 -1364
rect 6986 -1398 7020 -1364
rect 6276 -1431 7020 -1398
rect 6276 -1432 6377 -1431
rect 6276 -1466 6310 -1432
rect 6344 -1466 6377 -1432
rect 6276 -1500 6377 -1466
rect 6919 -1432 7020 -1431
rect 6919 -1466 6952 -1432
rect 6986 -1466 7020 -1432
rect 6276 -1534 6310 -1500
rect 6344 -1534 6377 -1500
rect 6276 -1568 6377 -1534
rect 6276 -1602 6310 -1568
rect 6344 -1602 6377 -1568
rect 6276 -1802 6377 -1602
rect 6276 -1836 6310 -1802
rect 6344 -1836 6377 -1802
rect 6276 -1870 6377 -1836
rect 6276 -1904 6310 -1870
rect 6344 -1904 6377 -1870
rect 6276 -1938 6377 -1904
rect 6919 -1500 7020 -1466
rect 6919 -1534 6952 -1500
rect 6986 -1534 7020 -1500
rect 6919 -1568 7020 -1534
rect 6919 -1602 6952 -1568
rect 6986 -1602 7020 -1568
rect 6919 -1802 7020 -1602
rect 6919 -1836 6952 -1802
rect 6986 -1836 7020 -1802
rect 6919 -1870 7020 -1836
rect 6919 -1904 6952 -1870
rect 6986 -1904 7020 -1870
rect 6276 -1972 6310 -1938
rect 6344 -1972 6377 -1938
rect 6276 -1973 6377 -1972
rect 6919 -1938 7020 -1904
rect 6919 -1972 6952 -1938
rect 6986 -1972 7020 -1938
rect 6919 -1973 7020 -1972
rect 6276 -2006 7020 -1973
rect 6276 -2040 6310 -2006
rect 6344 -2040 6378 -2006
rect 6412 -2040 6446 -2006
rect 6480 -2040 6514 -2006
rect 6548 -2040 6748 -2006
rect 6782 -2040 6816 -2006
rect 6850 -2040 6884 -2006
rect 6918 -2040 6952 -2006
rect 6986 -2040 7020 -2006
rect 6276 -2074 7020 -2040
rect -1104 -2184 -360 -2150
rect -1104 -2218 -1070 -2184
rect -1036 -2218 -1002 -2184
rect -968 -2218 -934 -2184
rect -900 -2218 -866 -2184
rect -832 -2218 -632 -2184
rect -598 -2218 -564 -2184
rect -530 -2218 -496 -2184
rect -462 -2218 -428 -2184
rect -394 -2218 -360 -2184
rect -1104 -2251 -360 -2218
rect -1104 -2252 -1003 -2251
rect -1104 -2286 -1070 -2252
rect -1036 -2286 -1003 -2252
rect -1104 -2320 -1003 -2286
rect -461 -2252 -360 -2251
rect -461 -2286 -428 -2252
rect -394 -2286 -360 -2252
rect -1104 -2354 -1070 -2320
rect -1036 -2354 -1003 -2320
rect -1104 -2388 -1003 -2354
rect -1104 -2422 -1070 -2388
rect -1036 -2422 -1003 -2388
rect -1104 -2622 -1003 -2422
rect -1104 -2656 -1070 -2622
rect -1036 -2656 -1003 -2622
rect -1104 -2690 -1003 -2656
rect -1104 -2724 -1070 -2690
rect -1036 -2724 -1003 -2690
rect -1104 -2758 -1003 -2724
rect -461 -2320 -360 -2286
rect -461 -2354 -428 -2320
rect -394 -2354 -360 -2320
rect -461 -2388 -360 -2354
rect -461 -2422 -428 -2388
rect -394 -2422 -360 -2388
rect -461 -2622 -360 -2422
rect -461 -2656 -428 -2622
rect -394 -2656 -360 -2622
rect -461 -2690 -360 -2656
rect -461 -2724 -428 -2690
rect -394 -2724 -360 -2690
rect -1104 -2792 -1070 -2758
rect -1036 -2792 -1003 -2758
rect -1104 -2793 -1003 -2792
rect -461 -2758 -360 -2724
rect -461 -2792 -428 -2758
rect -394 -2792 -360 -2758
rect -461 -2793 -360 -2792
rect -1104 -2826 -360 -2793
rect -1104 -2860 -1070 -2826
rect -1036 -2860 -1002 -2826
rect -968 -2860 -934 -2826
rect -900 -2860 -866 -2826
rect -832 -2860 -632 -2826
rect -598 -2860 -564 -2826
rect -530 -2860 -496 -2826
rect -462 -2860 -428 -2826
rect -394 -2860 -360 -2826
rect -1104 -2894 -360 -2860
rect -284 -2184 460 -2150
rect -284 -2218 -250 -2184
rect -216 -2218 -182 -2184
rect -148 -2218 -114 -2184
rect -80 -2218 -46 -2184
rect -12 -2218 188 -2184
rect 222 -2218 256 -2184
rect 290 -2218 324 -2184
rect 358 -2218 392 -2184
rect 426 -2218 460 -2184
rect -284 -2251 460 -2218
rect -284 -2252 -183 -2251
rect -284 -2286 -250 -2252
rect -216 -2286 -183 -2252
rect -284 -2320 -183 -2286
rect 359 -2252 460 -2251
rect 359 -2286 392 -2252
rect 426 -2286 460 -2252
rect -284 -2354 -250 -2320
rect -216 -2354 -183 -2320
rect -284 -2388 -183 -2354
rect -284 -2422 -250 -2388
rect -216 -2422 -183 -2388
rect -284 -2622 -183 -2422
rect -284 -2656 -250 -2622
rect -216 -2656 -183 -2622
rect -284 -2690 -183 -2656
rect -284 -2724 -250 -2690
rect -216 -2724 -183 -2690
rect -284 -2758 -183 -2724
rect 359 -2320 460 -2286
rect 359 -2354 392 -2320
rect 426 -2354 460 -2320
rect 359 -2388 460 -2354
rect 359 -2422 392 -2388
rect 426 -2422 460 -2388
rect 359 -2622 460 -2422
rect 359 -2656 392 -2622
rect 426 -2656 460 -2622
rect 359 -2690 460 -2656
rect 359 -2724 392 -2690
rect 426 -2724 460 -2690
rect -284 -2792 -250 -2758
rect -216 -2792 -183 -2758
rect -284 -2793 -183 -2792
rect 359 -2758 460 -2724
rect 359 -2792 392 -2758
rect 426 -2792 460 -2758
rect 359 -2793 460 -2792
rect -284 -2826 460 -2793
rect -284 -2860 -250 -2826
rect -216 -2860 -182 -2826
rect -148 -2860 -114 -2826
rect -80 -2860 -46 -2826
rect -12 -2860 188 -2826
rect 222 -2860 256 -2826
rect 290 -2860 324 -2826
rect 358 -2860 392 -2826
rect 426 -2860 460 -2826
rect -284 -2894 460 -2860
rect 536 -2184 1280 -2150
rect 536 -2218 570 -2184
rect 604 -2218 638 -2184
rect 672 -2218 706 -2184
rect 740 -2218 774 -2184
rect 808 -2218 1008 -2184
rect 1042 -2218 1076 -2184
rect 1110 -2218 1144 -2184
rect 1178 -2218 1212 -2184
rect 1246 -2218 1280 -2184
rect 536 -2251 1280 -2218
rect 536 -2252 637 -2251
rect 536 -2286 570 -2252
rect 604 -2286 637 -2252
rect 536 -2320 637 -2286
rect 1179 -2252 1280 -2251
rect 1179 -2286 1212 -2252
rect 1246 -2286 1280 -2252
rect 536 -2354 570 -2320
rect 604 -2354 637 -2320
rect 536 -2388 637 -2354
rect 536 -2422 570 -2388
rect 604 -2422 637 -2388
rect 536 -2622 637 -2422
rect 536 -2656 570 -2622
rect 604 -2656 637 -2622
rect 536 -2690 637 -2656
rect 536 -2724 570 -2690
rect 604 -2724 637 -2690
rect 536 -2758 637 -2724
rect 1179 -2320 1280 -2286
rect 1179 -2354 1212 -2320
rect 1246 -2354 1280 -2320
rect 1179 -2388 1280 -2354
rect 1179 -2422 1212 -2388
rect 1246 -2422 1280 -2388
rect 1179 -2622 1280 -2422
rect 1179 -2656 1212 -2622
rect 1246 -2656 1280 -2622
rect 1179 -2690 1280 -2656
rect 1179 -2724 1212 -2690
rect 1246 -2724 1280 -2690
rect 536 -2792 570 -2758
rect 604 -2792 637 -2758
rect 536 -2793 637 -2792
rect 1179 -2758 1280 -2724
rect 1179 -2792 1212 -2758
rect 1246 -2792 1280 -2758
rect 1179 -2793 1280 -2792
rect 536 -2826 1280 -2793
rect 536 -2860 570 -2826
rect 604 -2860 638 -2826
rect 672 -2860 706 -2826
rect 740 -2860 774 -2826
rect 808 -2860 1008 -2826
rect 1042 -2860 1076 -2826
rect 1110 -2860 1144 -2826
rect 1178 -2860 1212 -2826
rect 1246 -2860 1280 -2826
rect 536 -2894 1280 -2860
rect 1356 -2184 2100 -2150
rect 1356 -2218 1390 -2184
rect 1424 -2218 1458 -2184
rect 1492 -2218 1526 -2184
rect 1560 -2218 1594 -2184
rect 1628 -2218 1828 -2184
rect 1862 -2218 1896 -2184
rect 1930 -2218 1964 -2184
rect 1998 -2218 2032 -2184
rect 2066 -2218 2100 -2184
rect 1356 -2251 2100 -2218
rect 1356 -2252 1457 -2251
rect 1356 -2286 1390 -2252
rect 1424 -2286 1457 -2252
rect 1356 -2320 1457 -2286
rect 1999 -2252 2100 -2251
rect 1999 -2286 2032 -2252
rect 2066 -2286 2100 -2252
rect 1356 -2354 1390 -2320
rect 1424 -2354 1457 -2320
rect 1356 -2388 1457 -2354
rect 1356 -2422 1390 -2388
rect 1424 -2422 1457 -2388
rect 1356 -2622 1457 -2422
rect 1356 -2656 1390 -2622
rect 1424 -2656 1457 -2622
rect 1356 -2690 1457 -2656
rect 1356 -2724 1390 -2690
rect 1424 -2724 1457 -2690
rect 1356 -2758 1457 -2724
rect 1999 -2320 2100 -2286
rect 1999 -2354 2032 -2320
rect 2066 -2354 2100 -2320
rect 1999 -2388 2100 -2354
rect 1999 -2422 2032 -2388
rect 2066 -2422 2100 -2388
rect 1999 -2622 2100 -2422
rect 1999 -2656 2032 -2622
rect 2066 -2656 2100 -2622
rect 1999 -2690 2100 -2656
rect 1999 -2724 2032 -2690
rect 2066 -2724 2100 -2690
rect 1356 -2792 1390 -2758
rect 1424 -2792 1457 -2758
rect 1356 -2793 1457 -2792
rect 1999 -2758 2100 -2724
rect 1999 -2792 2032 -2758
rect 2066 -2792 2100 -2758
rect 1999 -2793 2100 -2792
rect 1356 -2826 2100 -2793
rect 1356 -2860 1390 -2826
rect 1424 -2860 1458 -2826
rect 1492 -2860 1526 -2826
rect 1560 -2860 1594 -2826
rect 1628 -2860 1828 -2826
rect 1862 -2860 1896 -2826
rect 1930 -2860 1964 -2826
rect 1998 -2860 2032 -2826
rect 2066 -2860 2100 -2826
rect 1356 -2894 2100 -2860
rect 2176 -2184 2920 -2150
rect 2176 -2218 2210 -2184
rect 2244 -2218 2278 -2184
rect 2312 -2218 2346 -2184
rect 2380 -2218 2414 -2184
rect 2448 -2218 2648 -2184
rect 2682 -2218 2716 -2184
rect 2750 -2218 2784 -2184
rect 2818 -2218 2852 -2184
rect 2886 -2218 2920 -2184
rect 2176 -2251 2920 -2218
rect 2176 -2252 2277 -2251
rect 2176 -2286 2210 -2252
rect 2244 -2286 2277 -2252
rect 2176 -2320 2277 -2286
rect 2819 -2252 2920 -2251
rect 2819 -2286 2852 -2252
rect 2886 -2286 2920 -2252
rect 2176 -2354 2210 -2320
rect 2244 -2354 2277 -2320
rect 2176 -2388 2277 -2354
rect 2176 -2422 2210 -2388
rect 2244 -2422 2277 -2388
rect 2176 -2622 2277 -2422
rect 2176 -2656 2210 -2622
rect 2244 -2656 2277 -2622
rect 2176 -2690 2277 -2656
rect 2176 -2724 2210 -2690
rect 2244 -2724 2277 -2690
rect 2176 -2758 2277 -2724
rect 2819 -2320 2920 -2286
rect 2819 -2354 2852 -2320
rect 2886 -2354 2920 -2320
rect 2819 -2388 2920 -2354
rect 2819 -2422 2852 -2388
rect 2886 -2422 2920 -2388
rect 2819 -2622 2920 -2422
rect 2819 -2656 2852 -2622
rect 2886 -2656 2920 -2622
rect 2819 -2690 2920 -2656
rect 2819 -2724 2852 -2690
rect 2886 -2724 2920 -2690
rect 2176 -2792 2210 -2758
rect 2244 -2792 2277 -2758
rect 2176 -2793 2277 -2792
rect 2819 -2758 2920 -2724
rect 2819 -2792 2852 -2758
rect 2886 -2792 2920 -2758
rect 2819 -2793 2920 -2792
rect 2176 -2826 2920 -2793
rect 2176 -2860 2210 -2826
rect 2244 -2860 2278 -2826
rect 2312 -2860 2346 -2826
rect 2380 -2860 2414 -2826
rect 2448 -2860 2648 -2826
rect 2682 -2860 2716 -2826
rect 2750 -2860 2784 -2826
rect 2818 -2860 2852 -2826
rect 2886 -2860 2920 -2826
rect 2176 -2894 2920 -2860
rect 2996 -2184 3740 -2150
rect 2996 -2218 3030 -2184
rect 3064 -2218 3098 -2184
rect 3132 -2218 3166 -2184
rect 3200 -2218 3234 -2184
rect 3268 -2218 3468 -2184
rect 3502 -2218 3536 -2184
rect 3570 -2218 3604 -2184
rect 3638 -2218 3672 -2184
rect 3706 -2218 3740 -2184
rect 2996 -2251 3740 -2218
rect 2996 -2252 3097 -2251
rect 2996 -2286 3030 -2252
rect 3064 -2286 3097 -2252
rect 2996 -2320 3097 -2286
rect 3639 -2252 3740 -2251
rect 3639 -2286 3672 -2252
rect 3706 -2286 3740 -2252
rect 2996 -2354 3030 -2320
rect 3064 -2354 3097 -2320
rect 2996 -2388 3097 -2354
rect 2996 -2422 3030 -2388
rect 3064 -2422 3097 -2388
rect 2996 -2622 3097 -2422
rect 2996 -2656 3030 -2622
rect 3064 -2656 3097 -2622
rect 2996 -2690 3097 -2656
rect 2996 -2724 3030 -2690
rect 3064 -2724 3097 -2690
rect 2996 -2758 3097 -2724
rect 3639 -2320 3740 -2286
rect 3639 -2354 3672 -2320
rect 3706 -2354 3740 -2320
rect 3639 -2388 3740 -2354
rect 3639 -2422 3672 -2388
rect 3706 -2422 3740 -2388
rect 3639 -2622 3740 -2422
rect 3639 -2656 3672 -2622
rect 3706 -2656 3740 -2622
rect 3639 -2690 3740 -2656
rect 3639 -2724 3672 -2690
rect 3706 -2724 3740 -2690
rect 2996 -2792 3030 -2758
rect 3064 -2792 3097 -2758
rect 2996 -2793 3097 -2792
rect 3639 -2758 3740 -2724
rect 3639 -2792 3672 -2758
rect 3706 -2792 3740 -2758
rect 3639 -2793 3740 -2792
rect 2996 -2826 3740 -2793
rect 2996 -2860 3030 -2826
rect 3064 -2860 3098 -2826
rect 3132 -2860 3166 -2826
rect 3200 -2860 3234 -2826
rect 3268 -2860 3468 -2826
rect 3502 -2860 3536 -2826
rect 3570 -2860 3604 -2826
rect 3638 -2860 3672 -2826
rect 3706 -2860 3740 -2826
rect 2996 -2894 3740 -2860
rect 3816 -2184 4560 -2150
rect 3816 -2218 3850 -2184
rect 3884 -2218 3918 -2184
rect 3952 -2218 3986 -2184
rect 4020 -2218 4054 -2184
rect 4088 -2218 4288 -2184
rect 4322 -2218 4356 -2184
rect 4390 -2218 4424 -2184
rect 4458 -2218 4492 -2184
rect 4526 -2218 4560 -2184
rect 3816 -2251 4560 -2218
rect 3816 -2252 3917 -2251
rect 3816 -2286 3850 -2252
rect 3884 -2286 3917 -2252
rect 3816 -2320 3917 -2286
rect 4459 -2252 4560 -2251
rect 4459 -2286 4492 -2252
rect 4526 -2286 4560 -2252
rect 3816 -2354 3850 -2320
rect 3884 -2354 3917 -2320
rect 3816 -2388 3917 -2354
rect 3816 -2422 3850 -2388
rect 3884 -2422 3917 -2388
rect 3816 -2622 3917 -2422
rect 3816 -2656 3850 -2622
rect 3884 -2656 3917 -2622
rect 3816 -2690 3917 -2656
rect 3816 -2724 3850 -2690
rect 3884 -2724 3917 -2690
rect 3816 -2758 3917 -2724
rect 4459 -2320 4560 -2286
rect 4459 -2354 4492 -2320
rect 4526 -2354 4560 -2320
rect 4459 -2388 4560 -2354
rect 4459 -2422 4492 -2388
rect 4526 -2422 4560 -2388
rect 4459 -2622 4560 -2422
rect 4459 -2656 4492 -2622
rect 4526 -2656 4560 -2622
rect 4459 -2690 4560 -2656
rect 4459 -2724 4492 -2690
rect 4526 -2724 4560 -2690
rect 3816 -2792 3850 -2758
rect 3884 -2792 3917 -2758
rect 3816 -2793 3917 -2792
rect 4459 -2758 4560 -2724
rect 4459 -2792 4492 -2758
rect 4526 -2792 4560 -2758
rect 4459 -2793 4560 -2792
rect 3816 -2826 4560 -2793
rect 3816 -2860 3850 -2826
rect 3884 -2860 3918 -2826
rect 3952 -2860 3986 -2826
rect 4020 -2860 4054 -2826
rect 4088 -2860 4288 -2826
rect 4322 -2860 4356 -2826
rect 4390 -2860 4424 -2826
rect 4458 -2860 4492 -2826
rect 4526 -2860 4560 -2826
rect 3816 -2894 4560 -2860
rect 4636 -2184 5380 -2150
rect 4636 -2218 4670 -2184
rect 4704 -2218 4738 -2184
rect 4772 -2218 4806 -2184
rect 4840 -2218 4874 -2184
rect 4908 -2218 5108 -2184
rect 5142 -2218 5176 -2184
rect 5210 -2218 5244 -2184
rect 5278 -2218 5312 -2184
rect 5346 -2218 5380 -2184
rect 4636 -2251 5380 -2218
rect 4636 -2252 4737 -2251
rect 4636 -2286 4670 -2252
rect 4704 -2286 4737 -2252
rect 4636 -2320 4737 -2286
rect 5279 -2252 5380 -2251
rect 5279 -2286 5312 -2252
rect 5346 -2286 5380 -2252
rect 4636 -2354 4670 -2320
rect 4704 -2354 4737 -2320
rect 4636 -2388 4737 -2354
rect 4636 -2422 4670 -2388
rect 4704 -2422 4737 -2388
rect 4636 -2622 4737 -2422
rect 4636 -2656 4670 -2622
rect 4704 -2656 4737 -2622
rect 4636 -2690 4737 -2656
rect 4636 -2724 4670 -2690
rect 4704 -2724 4737 -2690
rect 4636 -2758 4737 -2724
rect 5279 -2320 5380 -2286
rect 5279 -2354 5312 -2320
rect 5346 -2354 5380 -2320
rect 5279 -2388 5380 -2354
rect 5279 -2422 5312 -2388
rect 5346 -2422 5380 -2388
rect 5279 -2622 5380 -2422
rect 5279 -2656 5312 -2622
rect 5346 -2656 5380 -2622
rect 5279 -2690 5380 -2656
rect 5279 -2724 5312 -2690
rect 5346 -2724 5380 -2690
rect 4636 -2792 4670 -2758
rect 4704 -2792 4737 -2758
rect 4636 -2793 4737 -2792
rect 5279 -2758 5380 -2724
rect 5279 -2792 5312 -2758
rect 5346 -2792 5380 -2758
rect 5279 -2793 5380 -2792
rect 4636 -2826 5380 -2793
rect 4636 -2860 4670 -2826
rect 4704 -2860 4738 -2826
rect 4772 -2860 4806 -2826
rect 4840 -2860 4874 -2826
rect 4908 -2860 5108 -2826
rect 5142 -2860 5176 -2826
rect 5210 -2860 5244 -2826
rect 5278 -2860 5312 -2826
rect 5346 -2860 5380 -2826
rect 4636 -2894 5380 -2860
rect 5456 -2184 6200 -2150
rect 5456 -2218 5490 -2184
rect 5524 -2218 5558 -2184
rect 5592 -2218 5626 -2184
rect 5660 -2218 5694 -2184
rect 5728 -2218 5928 -2184
rect 5962 -2218 5996 -2184
rect 6030 -2218 6064 -2184
rect 6098 -2218 6132 -2184
rect 6166 -2218 6200 -2184
rect 5456 -2251 6200 -2218
rect 5456 -2252 5557 -2251
rect 5456 -2286 5490 -2252
rect 5524 -2286 5557 -2252
rect 5456 -2320 5557 -2286
rect 6099 -2252 6200 -2251
rect 6099 -2286 6132 -2252
rect 6166 -2286 6200 -2252
rect 5456 -2354 5490 -2320
rect 5524 -2354 5557 -2320
rect 5456 -2388 5557 -2354
rect 5456 -2422 5490 -2388
rect 5524 -2422 5557 -2388
rect 5456 -2622 5557 -2422
rect 5456 -2656 5490 -2622
rect 5524 -2656 5557 -2622
rect 5456 -2690 5557 -2656
rect 5456 -2724 5490 -2690
rect 5524 -2724 5557 -2690
rect 5456 -2758 5557 -2724
rect 6099 -2320 6200 -2286
rect 6099 -2354 6132 -2320
rect 6166 -2354 6200 -2320
rect 6099 -2388 6200 -2354
rect 6099 -2422 6132 -2388
rect 6166 -2422 6200 -2388
rect 6099 -2622 6200 -2422
rect 6099 -2656 6132 -2622
rect 6166 -2656 6200 -2622
rect 6099 -2690 6200 -2656
rect 6099 -2724 6132 -2690
rect 6166 -2724 6200 -2690
rect 5456 -2792 5490 -2758
rect 5524 -2792 5557 -2758
rect 5456 -2793 5557 -2792
rect 6099 -2758 6200 -2724
rect 6099 -2792 6132 -2758
rect 6166 -2792 6200 -2758
rect 6099 -2793 6200 -2792
rect 5456 -2826 6200 -2793
rect 5456 -2860 5490 -2826
rect 5524 -2860 5558 -2826
rect 5592 -2860 5626 -2826
rect 5660 -2860 5694 -2826
rect 5728 -2860 5928 -2826
rect 5962 -2860 5996 -2826
rect 6030 -2860 6064 -2826
rect 6098 -2860 6132 -2826
rect 6166 -2860 6200 -2826
rect 5456 -2894 6200 -2860
rect 6276 -2184 7020 -2150
rect 6276 -2218 6310 -2184
rect 6344 -2218 6378 -2184
rect 6412 -2218 6446 -2184
rect 6480 -2218 6514 -2184
rect 6548 -2218 6748 -2184
rect 6782 -2218 6816 -2184
rect 6850 -2218 6884 -2184
rect 6918 -2218 6952 -2184
rect 6986 -2218 7020 -2184
rect 6276 -2251 7020 -2218
rect 6276 -2252 6377 -2251
rect 6276 -2286 6310 -2252
rect 6344 -2286 6377 -2252
rect 6276 -2320 6377 -2286
rect 6919 -2252 7020 -2251
rect 6919 -2286 6952 -2252
rect 6986 -2286 7020 -2252
rect 6276 -2354 6310 -2320
rect 6344 -2354 6377 -2320
rect 6276 -2388 6377 -2354
rect 6276 -2422 6310 -2388
rect 6344 -2422 6377 -2388
rect 6276 -2622 6377 -2422
rect 6276 -2656 6310 -2622
rect 6344 -2656 6377 -2622
rect 6276 -2690 6377 -2656
rect 6276 -2724 6310 -2690
rect 6344 -2724 6377 -2690
rect 6276 -2758 6377 -2724
rect 6919 -2320 7020 -2286
rect 6919 -2354 6952 -2320
rect 6986 -2354 7020 -2320
rect 6919 -2388 7020 -2354
rect 6919 -2422 6952 -2388
rect 6986 -2422 7020 -2388
rect 6919 -2622 7020 -2422
rect 6919 -2656 6952 -2622
rect 6986 -2656 7020 -2622
rect 6919 -2690 7020 -2656
rect 6919 -2724 6952 -2690
rect 6986 -2724 7020 -2690
rect 6276 -2792 6310 -2758
rect 6344 -2792 6377 -2758
rect 6276 -2793 6377 -2792
rect 6919 -2758 7020 -2724
rect 6919 -2792 6952 -2758
rect 6986 -2792 7020 -2758
rect 6919 -2793 7020 -2792
rect 6276 -2826 7020 -2793
rect 6276 -2860 6310 -2826
rect 6344 -2860 6378 -2826
rect 6412 -2860 6446 -2826
rect 6480 -2860 6514 -2826
rect 6548 -2860 6748 -2826
rect 6782 -2860 6816 -2826
rect 6850 -2860 6884 -2826
rect 6918 -2860 6952 -2826
rect 6986 -2860 7020 -2826
rect 6276 -2894 7020 -2860
rect -1104 -3004 -360 -2970
rect -1104 -3038 -1070 -3004
rect -1036 -3038 -1002 -3004
rect -968 -3038 -934 -3004
rect -900 -3038 -866 -3004
rect -832 -3038 -632 -3004
rect -598 -3038 -564 -3004
rect -530 -3038 -496 -3004
rect -462 -3038 -428 -3004
rect -394 -3038 -360 -3004
rect -1104 -3071 -360 -3038
rect -1104 -3072 -1003 -3071
rect -1104 -3106 -1070 -3072
rect -1036 -3106 -1003 -3072
rect -1104 -3140 -1003 -3106
rect -461 -3072 -360 -3071
rect -461 -3106 -428 -3072
rect -394 -3106 -360 -3072
rect -1104 -3174 -1070 -3140
rect -1036 -3174 -1003 -3140
rect -1104 -3208 -1003 -3174
rect -1104 -3242 -1070 -3208
rect -1036 -3242 -1003 -3208
rect -1104 -3442 -1003 -3242
rect -1104 -3476 -1070 -3442
rect -1036 -3476 -1003 -3442
rect -1104 -3510 -1003 -3476
rect -1104 -3544 -1070 -3510
rect -1036 -3544 -1003 -3510
rect -1104 -3578 -1003 -3544
rect -461 -3140 -360 -3106
rect -461 -3174 -428 -3140
rect -394 -3174 -360 -3140
rect -461 -3208 -360 -3174
rect -461 -3242 -428 -3208
rect -394 -3242 -360 -3208
rect -461 -3442 -360 -3242
rect -461 -3476 -428 -3442
rect -394 -3476 -360 -3442
rect -461 -3510 -360 -3476
rect -461 -3544 -428 -3510
rect -394 -3544 -360 -3510
rect -1104 -3612 -1070 -3578
rect -1036 -3612 -1003 -3578
rect -1104 -3613 -1003 -3612
rect -461 -3578 -360 -3544
rect -461 -3612 -428 -3578
rect -394 -3612 -360 -3578
rect -461 -3613 -360 -3612
rect -1104 -3646 -360 -3613
rect -1104 -3680 -1070 -3646
rect -1036 -3680 -1002 -3646
rect -968 -3680 -934 -3646
rect -900 -3680 -866 -3646
rect -832 -3680 -632 -3646
rect -598 -3680 -564 -3646
rect -530 -3680 -496 -3646
rect -462 -3680 -428 -3646
rect -394 -3680 -360 -3646
rect -1104 -3714 -360 -3680
rect -284 -3004 460 -2970
rect -284 -3038 -250 -3004
rect -216 -3038 -182 -3004
rect -148 -3038 -114 -3004
rect -80 -3038 -46 -3004
rect -12 -3038 188 -3004
rect 222 -3038 256 -3004
rect 290 -3038 324 -3004
rect 358 -3038 392 -3004
rect 426 -3038 460 -3004
rect -284 -3071 460 -3038
rect -284 -3072 -183 -3071
rect -284 -3106 -250 -3072
rect -216 -3106 -183 -3072
rect -284 -3140 -183 -3106
rect 359 -3072 460 -3071
rect 359 -3106 392 -3072
rect 426 -3106 460 -3072
rect -284 -3174 -250 -3140
rect -216 -3174 -183 -3140
rect -284 -3208 -183 -3174
rect -284 -3242 -250 -3208
rect -216 -3242 -183 -3208
rect -284 -3442 -183 -3242
rect -284 -3476 -250 -3442
rect -216 -3476 -183 -3442
rect -284 -3510 -183 -3476
rect -284 -3544 -250 -3510
rect -216 -3544 -183 -3510
rect -284 -3578 -183 -3544
rect 359 -3140 460 -3106
rect 359 -3174 392 -3140
rect 426 -3174 460 -3140
rect 359 -3208 460 -3174
rect 359 -3242 392 -3208
rect 426 -3242 460 -3208
rect 359 -3442 460 -3242
rect 359 -3476 392 -3442
rect 426 -3476 460 -3442
rect 359 -3510 460 -3476
rect 359 -3544 392 -3510
rect 426 -3544 460 -3510
rect -284 -3612 -250 -3578
rect -216 -3612 -183 -3578
rect -284 -3613 -183 -3612
rect 359 -3578 460 -3544
rect 359 -3612 392 -3578
rect 426 -3612 460 -3578
rect 359 -3613 460 -3612
rect -284 -3646 460 -3613
rect -284 -3680 -250 -3646
rect -216 -3680 -182 -3646
rect -148 -3680 -114 -3646
rect -80 -3680 -46 -3646
rect -12 -3680 188 -3646
rect 222 -3680 256 -3646
rect 290 -3680 324 -3646
rect 358 -3680 392 -3646
rect 426 -3680 460 -3646
rect -284 -3714 460 -3680
rect 536 -3004 1280 -2970
rect 536 -3038 570 -3004
rect 604 -3038 638 -3004
rect 672 -3038 706 -3004
rect 740 -3038 774 -3004
rect 808 -3038 1008 -3004
rect 1042 -3038 1076 -3004
rect 1110 -3038 1144 -3004
rect 1178 -3038 1212 -3004
rect 1246 -3038 1280 -3004
rect 536 -3071 1280 -3038
rect 536 -3072 637 -3071
rect 536 -3106 570 -3072
rect 604 -3106 637 -3072
rect 536 -3140 637 -3106
rect 1179 -3072 1280 -3071
rect 1179 -3106 1212 -3072
rect 1246 -3106 1280 -3072
rect 536 -3174 570 -3140
rect 604 -3174 637 -3140
rect 536 -3208 637 -3174
rect 536 -3242 570 -3208
rect 604 -3242 637 -3208
rect 536 -3442 637 -3242
rect 536 -3476 570 -3442
rect 604 -3476 637 -3442
rect 536 -3510 637 -3476
rect 536 -3544 570 -3510
rect 604 -3544 637 -3510
rect 536 -3578 637 -3544
rect 1179 -3140 1280 -3106
rect 1179 -3174 1212 -3140
rect 1246 -3174 1280 -3140
rect 1179 -3208 1280 -3174
rect 1179 -3242 1212 -3208
rect 1246 -3242 1280 -3208
rect 1179 -3442 1280 -3242
rect 1179 -3476 1212 -3442
rect 1246 -3476 1280 -3442
rect 1179 -3510 1280 -3476
rect 1179 -3544 1212 -3510
rect 1246 -3544 1280 -3510
rect 536 -3612 570 -3578
rect 604 -3612 637 -3578
rect 536 -3613 637 -3612
rect 1179 -3578 1280 -3544
rect 1179 -3612 1212 -3578
rect 1246 -3612 1280 -3578
rect 1179 -3613 1280 -3612
rect 536 -3646 1280 -3613
rect 536 -3680 570 -3646
rect 604 -3680 638 -3646
rect 672 -3680 706 -3646
rect 740 -3680 774 -3646
rect 808 -3680 1008 -3646
rect 1042 -3680 1076 -3646
rect 1110 -3680 1144 -3646
rect 1178 -3680 1212 -3646
rect 1246 -3680 1280 -3646
rect 536 -3714 1280 -3680
rect 1356 -3004 2100 -2970
rect 1356 -3038 1390 -3004
rect 1424 -3038 1458 -3004
rect 1492 -3038 1526 -3004
rect 1560 -3038 1594 -3004
rect 1628 -3038 1828 -3004
rect 1862 -3038 1896 -3004
rect 1930 -3038 1964 -3004
rect 1998 -3038 2032 -3004
rect 2066 -3038 2100 -3004
rect 1356 -3071 2100 -3038
rect 1356 -3072 1457 -3071
rect 1356 -3106 1390 -3072
rect 1424 -3106 1457 -3072
rect 1356 -3140 1457 -3106
rect 1999 -3072 2100 -3071
rect 1999 -3106 2032 -3072
rect 2066 -3106 2100 -3072
rect 1356 -3174 1390 -3140
rect 1424 -3174 1457 -3140
rect 1356 -3208 1457 -3174
rect 1356 -3242 1390 -3208
rect 1424 -3242 1457 -3208
rect 1356 -3442 1457 -3242
rect 1356 -3476 1390 -3442
rect 1424 -3476 1457 -3442
rect 1356 -3510 1457 -3476
rect 1356 -3544 1390 -3510
rect 1424 -3544 1457 -3510
rect 1356 -3578 1457 -3544
rect 1999 -3140 2100 -3106
rect 1999 -3174 2032 -3140
rect 2066 -3174 2100 -3140
rect 1999 -3208 2100 -3174
rect 1999 -3242 2032 -3208
rect 2066 -3242 2100 -3208
rect 1999 -3442 2100 -3242
rect 1999 -3476 2032 -3442
rect 2066 -3476 2100 -3442
rect 1999 -3510 2100 -3476
rect 1999 -3544 2032 -3510
rect 2066 -3544 2100 -3510
rect 1356 -3612 1390 -3578
rect 1424 -3612 1457 -3578
rect 1356 -3613 1457 -3612
rect 1999 -3578 2100 -3544
rect 1999 -3612 2032 -3578
rect 2066 -3612 2100 -3578
rect 1999 -3613 2100 -3612
rect 1356 -3646 2100 -3613
rect 1356 -3680 1390 -3646
rect 1424 -3680 1458 -3646
rect 1492 -3680 1526 -3646
rect 1560 -3680 1594 -3646
rect 1628 -3680 1828 -3646
rect 1862 -3680 1896 -3646
rect 1930 -3680 1964 -3646
rect 1998 -3680 2032 -3646
rect 2066 -3680 2100 -3646
rect 1356 -3714 2100 -3680
rect 2176 -3004 2920 -2970
rect 2176 -3038 2210 -3004
rect 2244 -3038 2278 -3004
rect 2312 -3038 2346 -3004
rect 2380 -3038 2414 -3004
rect 2448 -3038 2648 -3004
rect 2682 -3038 2716 -3004
rect 2750 -3038 2784 -3004
rect 2818 -3038 2852 -3004
rect 2886 -3038 2920 -3004
rect 2176 -3071 2920 -3038
rect 2176 -3072 2277 -3071
rect 2176 -3106 2210 -3072
rect 2244 -3106 2277 -3072
rect 2176 -3140 2277 -3106
rect 2819 -3072 2920 -3071
rect 2819 -3106 2852 -3072
rect 2886 -3106 2920 -3072
rect 2176 -3174 2210 -3140
rect 2244 -3174 2277 -3140
rect 2176 -3208 2277 -3174
rect 2176 -3242 2210 -3208
rect 2244 -3242 2277 -3208
rect 2176 -3442 2277 -3242
rect 2176 -3476 2210 -3442
rect 2244 -3476 2277 -3442
rect 2176 -3510 2277 -3476
rect 2176 -3544 2210 -3510
rect 2244 -3544 2277 -3510
rect 2176 -3578 2277 -3544
rect 2819 -3140 2920 -3106
rect 2819 -3174 2852 -3140
rect 2886 -3174 2920 -3140
rect 2819 -3208 2920 -3174
rect 2819 -3242 2852 -3208
rect 2886 -3242 2920 -3208
rect 2819 -3442 2920 -3242
rect 2819 -3476 2852 -3442
rect 2886 -3476 2920 -3442
rect 2819 -3510 2920 -3476
rect 2819 -3544 2852 -3510
rect 2886 -3544 2920 -3510
rect 2176 -3612 2210 -3578
rect 2244 -3612 2277 -3578
rect 2176 -3613 2277 -3612
rect 2819 -3578 2920 -3544
rect 2819 -3612 2852 -3578
rect 2886 -3612 2920 -3578
rect 2819 -3613 2920 -3612
rect 2176 -3646 2920 -3613
rect 2176 -3680 2210 -3646
rect 2244 -3680 2278 -3646
rect 2312 -3680 2346 -3646
rect 2380 -3680 2414 -3646
rect 2448 -3680 2648 -3646
rect 2682 -3680 2716 -3646
rect 2750 -3680 2784 -3646
rect 2818 -3680 2852 -3646
rect 2886 -3680 2920 -3646
rect 2176 -3714 2920 -3680
rect 2996 -3004 3740 -2970
rect 2996 -3038 3030 -3004
rect 3064 -3038 3098 -3004
rect 3132 -3038 3166 -3004
rect 3200 -3038 3234 -3004
rect 3268 -3038 3468 -3004
rect 3502 -3038 3536 -3004
rect 3570 -3038 3604 -3004
rect 3638 -3038 3672 -3004
rect 3706 -3038 3740 -3004
rect 2996 -3071 3740 -3038
rect 2996 -3072 3097 -3071
rect 2996 -3106 3030 -3072
rect 3064 -3106 3097 -3072
rect 2996 -3140 3097 -3106
rect 3639 -3072 3740 -3071
rect 3639 -3106 3672 -3072
rect 3706 -3106 3740 -3072
rect 2996 -3174 3030 -3140
rect 3064 -3174 3097 -3140
rect 2996 -3208 3097 -3174
rect 2996 -3242 3030 -3208
rect 3064 -3242 3097 -3208
rect 2996 -3442 3097 -3242
rect 2996 -3476 3030 -3442
rect 3064 -3476 3097 -3442
rect 2996 -3510 3097 -3476
rect 2996 -3544 3030 -3510
rect 3064 -3544 3097 -3510
rect 2996 -3578 3097 -3544
rect 3639 -3140 3740 -3106
rect 3639 -3174 3672 -3140
rect 3706 -3174 3740 -3140
rect 3639 -3208 3740 -3174
rect 3639 -3242 3672 -3208
rect 3706 -3242 3740 -3208
rect 3639 -3442 3740 -3242
rect 3639 -3476 3672 -3442
rect 3706 -3476 3740 -3442
rect 3639 -3510 3740 -3476
rect 3639 -3544 3672 -3510
rect 3706 -3544 3740 -3510
rect 2996 -3612 3030 -3578
rect 3064 -3612 3097 -3578
rect 2996 -3613 3097 -3612
rect 3639 -3578 3740 -3544
rect 3639 -3612 3672 -3578
rect 3706 -3612 3740 -3578
rect 3639 -3613 3740 -3612
rect 2996 -3646 3740 -3613
rect 2996 -3680 3030 -3646
rect 3064 -3680 3098 -3646
rect 3132 -3680 3166 -3646
rect 3200 -3680 3234 -3646
rect 3268 -3680 3468 -3646
rect 3502 -3680 3536 -3646
rect 3570 -3680 3604 -3646
rect 3638 -3680 3672 -3646
rect 3706 -3680 3740 -3646
rect 2996 -3714 3740 -3680
rect 3816 -3004 4560 -2970
rect 3816 -3038 3850 -3004
rect 3884 -3038 3918 -3004
rect 3952 -3038 3986 -3004
rect 4020 -3038 4054 -3004
rect 4088 -3038 4288 -3004
rect 4322 -3038 4356 -3004
rect 4390 -3038 4424 -3004
rect 4458 -3038 4492 -3004
rect 4526 -3038 4560 -3004
rect 3816 -3071 4560 -3038
rect 3816 -3072 3917 -3071
rect 3816 -3106 3850 -3072
rect 3884 -3106 3917 -3072
rect 3816 -3140 3917 -3106
rect 4459 -3072 4560 -3071
rect 4459 -3106 4492 -3072
rect 4526 -3106 4560 -3072
rect 3816 -3174 3850 -3140
rect 3884 -3174 3917 -3140
rect 3816 -3208 3917 -3174
rect 3816 -3242 3850 -3208
rect 3884 -3242 3917 -3208
rect 3816 -3442 3917 -3242
rect 3816 -3476 3850 -3442
rect 3884 -3476 3917 -3442
rect 3816 -3510 3917 -3476
rect 3816 -3544 3850 -3510
rect 3884 -3544 3917 -3510
rect 3816 -3578 3917 -3544
rect 4459 -3140 4560 -3106
rect 4459 -3174 4492 -3140
rect 4526 -3174 4560 -3140
rect 4459 -3208 4560 -3174
rect 4459 -3242 4492 -3208
rect 4526 -3242 4560 -3208
rect 4459 -3442 4560 -3242
rect 4459 -3476 4492 -3442
rect 4526 -3476 4560 -3442
rect 4459 -3510 4560 -3476
rect 4459 -3544 4492 -3510
rect 4526 -3544 4560 -3510
rect 3816 -3612 3850 -3578
rect 3884 -3612 3917 -3578
rect 3816 -3613 3917 -3612
rect 4459 -3578 4560 -3544
rect 4459 -3612 4492 -3578
rect 4526 -3612 4560 -3578
rect 4459 -3613 4560 -3612
rect 3816 -3646 4560 -3613
rect 3816 -3680 3850 -3646
rect 3884 -3680 3918 -3646
rect 3952 -3680 3986 -3646
rect 4020 -3680 4054 -3646
rect 4088 -3680 4288 -3646
rect 4322 -3680 4356 -3646
rect 4390 -3680 4424 -3646
rect 4458 -3680 4492 -3646
rect 4526 -3680 4560 -3646
rect 3816 -3714 4560 -3680
rect 4636 -3004 5380 -2970
rect 4636 -3038 4670 -3004
rect 4704 -3038 4738 -3004
rect 4772 -3038 4806 -3004
rect 4840 -3038 4874 -3004
rect 4908 -3038 5108 -3004
rect 5142 -3038 5176 -3004
rect 5210 -3038 5244 -3004
rect 5278 -3038 5312 -3004
rect 5346 -3038 5380 -3004
rect 4636 -3071 5380 -3038
rect 4636 -3072 4737 -3071
rect 4636 -3106 4670 -3072
rect 4704 -3106 4737 -3072
rect 4636 -3140 4737 -3106
rect 5279 -3072 5380 -3071
rect 5279 -3106 5312 -3072
rect 5346 -3106 5380 -3072
rect 4636 -3174 4670 -3140
rect 4704 -3174 4737 -3140
rect 4636 -3208 4737 -3174
rect 4636 -3242 4670 -3208
rect 4704 -3242 4737 -3208
rect 4636 -3442 4737 -3242
rect 4636 -3476 4670 -3442
rect 4704 -3476 4737 -3442
rect 4636 -3510 4737 -3476
rect 4636 -3544 4670 -3510
rect 4704 -3544 4737 -3510
rect 4636 -3578 4737 -3544
rect 5279 -3140 5380 -3106
rect 5279 -3174 5312 -3140
rect 5346 -3174 5380 -3140
rect 5279 -3208 5380 -3174
rect 5279 -3242 5312 -3208
rect 5346 -3242 5380 -3208
rect 5279 -3442 5380 -3242
rect 5279 -3476 5312 -3442
rect 5346 -3476 5380 -3442
rect 5279 -3510 5380 -3476
rect 5279 -3544 5312 -3510
rect 5346 -3544 5380 -3510
rect 4636 -3612 4670 -3578
rect 4704 -3612 4737 -3578
rect 4636 -3613 4737 -3612
rect 5279 -3578 5380 -3544
rect 5279 -3612 5312 -3578
rect 5346 -3612 5380 -3578
rect 5279 -3613 5380 -3612
rect 4636 -3646 5380 -3613
rect 4636 -3680 4670 -3646
rect 4704 -3680 4738 -3646
rect 4772 -3680 4806 -3646
rect 4840 -3680 4874 -3646
rect 4908 -3680 5108 -3646
rect 5142 -3680 5176 -3646
rect 5210 -3680 5244 -3646
rect 5278 -3680 5312 -3646
rect 5346 -3680 5380 -3646
rect 4636 -3714 5380 -3680
rect 5456 -3004 6200 -2970
rect 5456 -3038 5490 -3004
rect 5524 -3038 5558 -3004
rect 5592 -3038 5626 -3004
rect 5660 -3038 5694 -3004
rect 5728 -3038 5928 -3004
rect 5962 -3038 5996 -3004
rect 6030 -3038 6064 -3004
rect 6098 -3038 6132 -3004
rect 6166 -3038 6200 -3004
rect 5456 -3071 6200 -3038
rect 5456 -3072 5557 -3071
rect 5456 -3106 5490 -3072
rect 5524 -3106 5557 -3072
rect 5456 -3140 5557 -3106
rect 6099 -3072 6200 -3071
rect 6099 -3106 6132 -3072
rect 6166 -3106 6200 -3072
rect 5456 -3174 5490 -3140
rect 5524 -3174 5557 -3140
rect 5456 -3208 5557 -3174
rect 5456 -3242 5490 -3208
rect 5524 -3242 5557 -3208
rect 5456 -3442 5557 -3242
rect 5456 -3476 5490 -3442
rect 5524 -3476 5557 -3442
rect 5456 -3510 5557 -3476
rect 5456 -3544 5490 -3510
rect 5524 -3544 5557 -3510
rect 5456 -3578 5557 -3544
rect 6099 -3140 6200 -3106
rect 6099 -3174 6132 -3140
rect 6166 -3174 6200 -3140
rect 6099 -3208 6200 -3174
rect 6099 -3242 6132 -3208
rect 6166 -3242 6200 -3208
rect 6099 -3442 6200 -3242
rect 6099 -3476 6132 -3442
rect 6166 -3476 6200 -3442
rect 6099 -3510 6200 -3476
rect 6099 -3544 6132 -3510
rect 6166 -3544 6200 -3510
rect 5456 -3612 5490 -3578
rect 5524 -3612 5557 -3578
rect 5456 -3613 5557 -3612
rect 6099 -3578 6200 -3544
rect 6099 -3612 6132 -3578
rect 6166 -3612 6200 -3578
rect 6099 -3613 6200 -3612
rect 5456 -3646 6200 -3613
rect 5456 -3680 5490 -3646
rect 5524 -3680 5558 -3646
rect 5592 -3680 5626 -3646
rect 5660 -3680 5694 -3646
rect 5728 -3680 5928 -3646
rect 5962 -3680 5996 -3646
rect 6030 -3680 6064 -3646
rect 6098 -3680 6132 -3646
rect 6166 -3680 6200 -3646
rect 5456 -3714 6200 -3680
rect 6276 -3004 7020 -2970
rect 6276 -3038 6310 -3004
rect 6344 -3038 6378 -3004
rect 6412 -3038 6446 -3004
rect 6480 -3038 6514 -3004
rect 6548 -3038 6748 -3004
rect 6782 -3038 6816 -3004
rect 6850 -3038 6884 -3004
rect 6918 -3038 6952 -3004
rect 6986 -3038 7020 -3004
rect 6276 -3071 7020 -3038
rect 6276 -3072 6377 -3071
rect 6276 -3106 6310 -3072
rect 6344 -3106 6377 -3072
rect 6276 -3140 6377 -3106
rect 6919 -3072 7020 -3071
rect 6919 -3106 6952 -3072
rect 6986 -3106 7020 -3072
rect 6276 -3174 6310 -3140
rect 6344 -3174 6377 -3140
rect 6276 -3208 6377 -3174
rect 6276 -3242 6310 -3208
rect 6344 -3242 6377 -3208
rect 6276 -3442 6377 -3242
rect 6276 -3476 6310 -3442
rect 6344 -3476 6377 -3442
rect 6276 -3510 6377 -3476
rect 6276 -3544 6310 -3510
rect 6344 -3544 6377 -3510
rect 6276 -3578 6377 -3544
rect 6919 -3140 7020 -3106
rect 6919 -3174 6952 -3140
rect 6986 -3174 7020 -3140
rect 6919 -3208 7020 -3174
rect 6919 -3242 6952 -3208
rect 6986 -3242 7020 -3208
rect 6919 -3442 7020 -3242
rect 6919 -3476 6952 -3442
rect 6986 -3476 7020 -3442
rect 6919 -3510 7020 -3476
rect 6919 -3544 6952 -3510
rect 6986 -3544 7020 -3510
rect 6276 -3612 6310 -3578
rect 6344 -3612 6377 -3578
rect 6276 -3613 6377 -3612
rect 6919 -3578 7020 -3544
rect 6919 -3612 6952 -3578
rect 6986 -3612 7020 -3578
rect 6919 -3613 7020 -3612
rect 6276 -3646 7020 -3613
rect 6276 -3680 6310 -3646
rect 6344 -3680 6378 -3646
rect 6412 -3680 6446 -3646
rect 6480 -3680 6514 -3646
rect 6548 -3680 6748 -3646
rect 6782 -3680 6816 -3646
rect 6850 -3680 6884 -3646
rect 6918 -3680 6952 -3646
rect 6986 -3680 7020 -3646
rect 6276 -3714 7020 -3680
rect -1104 -3824 -360 -3790
rect -1104 -3858 -1070 -3824
rect -1036 -3858 -1002 -3824
rect -968 -3858 -934 -3824
rect -900 -3858 -866 -3824
rect -832 -3858 -632 -3824
rect -598 -3858 -564 -3824
rect -530 -3858 -496 -3824
rect -462 -3858 -428 -3824
rect -394 -3858 -360 -3824
rect -1104 -3891 -360 -3858
rect -1104 -3892 -1003 -3891
rect -1104 -3926 -1070 -3892
rect -1036 -3926 -1003 -3892
rect -1104 -3960 -1003 -3926
rect -461 -3892 -360 -3891
rect -461 -3926 -428 -3892
rect -394 -3926 -360 -3892
rect -1104 -3994 -1070 -3960
rect -1036 -3994 -1003 -3960
rect -1104 -4028 -1003 -3994
rect -1104 -4062 -1070 -4028
rect -1036 -4062 -1003 -4028
rect -1104 -4262 -1003 -4062
rect -1104 -4296 -1070 -4262
rect -1036 -4296 -1003 -4262
rect -1104 -4330 -1003 -4296
rect -1104 -4364 -1070 -4330
rect -1036 -4364 -1003 -4330
rect -1104 -4398 -1003 -4364
rect -461 -3960 -360 -3926
rect -461 -3994 -428 -3960
rect -394 -3994 -360 -3960
rect -461 -4028 -360 -3994
rect -461 -4062 -428 -4028
rect -394 -4062 -360 -4028
rect -461 -4262 -360 -4062
rect -461 -4296 -428 -4262
rect -394 -4296 -360 -4262
rect -461 -4330 -360 -4296
rect -461 -4364 -428 -4330
rect -394 -4364 -360 -4330
rect -1104 -4432 -1070 -4398
rect -1036 -4432 -1003 -4398
rect -1104 -4433 -1003 -4432
rect -461 -4398 -360 -4364
rect -461 -4432 -428 -4398
rect -394 -4432 -360 -4398
rect -461 -4433 -360 -4432
rect -1104 -4466 -360 -4433
rect -1104 -4500 -1070 -4466
rect -1036 -4500 -1002 -4466
rect -968 -4500 -934 -4466
rect -900 -4500 -866 -4466
rect -832 -4500 -632 -4466
rect -598 -4500 -564 -4466
rect -530 -4500 -496 -4466
rect -462 -4500 -428 -4466
rect -394 -4500 -360 -4466
rect -1104 -4534 -360 -4500
rect -284 -3824 460 -3790
rect -284 -3858 -250 -3824
rect -216 -3858 -182 -3824
rect -148 -3858 -114 -3824
rect -80 -3858 -46 -3824
rect -12 -3858 188 -3824
rect 222 -3858 256 -3824
rect 290 -3858 324 -3824
rect 358 -3858 392 -3824
rect 426 -3858 460 -3824
rect -284 -3891 460 -3858
rect -284 -3892 -183 -3891
rect -284 -3926 -250 -3892
rect -216 -3926 -183 -3892
rect -284 -3960 -183 -3926
rect 359 -3892 460 -3891
rect 359 -3926 392 -3892
rect 426 -3926 460 -3892
rect -284 -3994 -250 -3960
rect -216 -3994 -183 -3960
rect -284 -4028 -183 -3994
rect -284 -4062 -250 -4028
rect -216 -4062 -183 -4028
rect -284 -4262 -183 -4062
rect -284 -4296 -250 -4262
rect -216 -4296 -183 -4262
rect -284 -4330 -183 -4296
rect -284 -4364 -250 -4330
rect -216 -4364 -183 -4330
rect -284 -4398 -183 -4364
rect 359 -3960 460 -3926
rect 359 -3994 392 -3960
rect 426 -3994 460 -3960
rect 359 -4028 460 -3994
rect 359 -4062 392 -4028
rect 426 -4062 460 -4028
rect 359 -4262 460 -4062
rect 359 -4296 392 -4262
rect 426 -4296 460 -4262
rect 359 -4330 460 -4296
rect 359 -4364 392 -4330
rect 426 -4364 460 -4330
rect -284 -4432 -250 -4398
rect -216 -4432 -183 -4398
rect -284 -4433 -183 -4432
rect 359 -4398 460 -4364
rect 359 -4432 392 -4398
rect 426 -4432 460 -4398
rect 359 -4433 460 -4432
rect -284 -4466 460 -4433
rect -284 -4500 -250 -4466
rect -216 -4500 -182 -4466
rect -148 -4500 -114 -4466
rect -80 -4500 -46 -4466
rect -12 -4500 188 -4466
rect 222 -4500 256 -4466
rect 290 -4500 324 -4466
rect 358 -4500 392 -4466
rect 426 -4500 460 -4466
rect -284 -4534 460 -4500
rect 536 -3824 1280 -3790
rect 536 -3858 570 -3824
rect 604 -3858 638 -3824
rect 672 -3858 706 -3824
rect 740 -3858 774 -3824
rect 808 -3858 1008 -3824
rect 1042 -3858 1076 -3824
rect 1110 -3858 1144 -3824
rect 1178 -3858 1212 -3824
rect 1246 -3858 1280 -3824
rect 536 -3891 1280 -3858
rect 536 -3892 637 -3891
rect 536 -3926 570 -3892
rect 604 -3926 637 -3892
rect 536 -3960 637 -3926
rect 1179 -3892 1280 -3891
rect 1179 -3926 1212 -3892
rect 1246 -3926 1280 -3892
rect 536 -3994 570 -3960
rect 604 -3994 637 -3960
rect 536 -4028 637 -3994
rect 536 -4062 570 -4028
rect 604 -4062 637 -4028
rect 536 -4262 637 -4062
rect 536 -4296 570 -4262
rect 604 -4296 637 -4262
rect 536 -4330 637 -4296
rect 536 -4364 570 -4330
rect 604 -4364 637 -4330
rect 536 -4398 637 -4364
rect 1179 -3960 1280 -3926
rect 1179 -3994 1212 -3960
rect 1246 -3994 1280 -3960
rect 1179 -4028 1280 -3994
rect 1179 -4062 1212 -4028
rect 1246 -4062 1280 -4028
rect 1179 -4262 1280 -4062
rect 1179 -4296 1212 -4262
rect 1246 -4296 1280 -4262
rect 1179 -4330 1280 -4296
rect 1179 -4364 1212 -4330
rect 1246 -4364 1280 -4330
rect 536 -4432 570 -4398
rect 604 -4432 637 -4398
rect 536 -4433 637 -4432
rect 1179 -4398 1280 -4364
rect 1179 -4432 1212 -4398
rect 1246 -4432 1280 -4398
rect 1179 -4433 1280 -4432
rect 536 -4466 1280 -4433
rect 536 -4500 570 -4466
rect 604 -4500 638 -4466
rect 672 -4500 706 -4466
rect 740 -4500 774 -4466
rect 808 -4500 1008 -4466
rect 1042 -4500 1076 -4466
rect 1110 -4500 1144 -4466
rect 1178 -4500 1212 -4466
rect 1246 -4500 1280 -4466
rect 536 -4534 1280 -4500
rect 1356 -3824 2100 -3790
rect 1356 -3858 1390 -3824
rect 1424 -3858 1458 -3824
rect 1492 -3858 1526 -3824
rect 1560 -3858 1594 -3824
rect 1628 -3858 1828 -3824
rect 1862 -3858 1896 -3824
rect 1930 -3858 1964 -3824
rect 1998 -3858 2032 -3824
rect 2066 -3858 2100 -3824
rect 1356 -3891 2100 -3858
rect 1356 -3892 1457 -3891
rect 1356 -3926 1390 -3892
rect 1424 -3926 1457 -3892
rect 1356 -3960 1457 -3926
rect 1999 -3892 2100 -3891
rect 1999 -3926 2032 -3892
rect 2066 -3926 2100 -3892
rect 1356 -3994 1390 -3960
rect 1424 -3994 1457 -3960
rect 1356 -4028 1457 -3994
rect 1356 -4062 1390 -4028
rect 1424 -4062 1457 -4028
rect 1356 -4262 1457 -4062
rect 1356 -4296 1390 -4262
rect 1424 -4296 1457 -4262
rect 1356 -4330 1457 -4296
rect 1356 -4364 1390 -4330
rect 1424 -4364 1457 -4330
rect 1356 -4398 1457 -4364
rect 1999 -3960 2100 -3926
rect 1999 -3994 2032 -3960
rect 2066 -3994 2100 -3960
rect 1999 -4028 2100 -3994
rect 1999 -4062 2032 -4028
rect 2066 -4062 2100 -4028
rect 1999 -4262 2100 -4062
rect 1999 -4296 2032 -4262
rect 2066 -4296 2100 -4262
rect 1999 -4330 2100 -4296
rect 1999 -4364 2032 -4330
rect 2066 -4364 2100 -4330
rect 1356 -4432 1390 -4398
rect 1424 -4432 1457 -4398
rect 1356 -4433 1457 -4432
rect 1999 -4398 2100 -4364
rect 1999 -4432 2032 -4398
rect 2066 -4432 2100 -4398
rect 1999 -4433 2100 -4432
rect 1356 -4466 2100 -4433
rect 1356 -4500 1390 -4466
rect 1424 -4500 1458 -4466
rect 1492 -4500 1526 -4466
rect 1560 -4500 1594 -4466
rect 1628 -4500 1828 -4466
rect 1862 -4500 1896 -4466
rect 1930 -4500 1964 -4466
rect 1998 -4500 2032 -4466
rect 2066 -4500 2100 -4466
rect 1356 -4534 2100 -4500
rect 2176 -3824 2920 -3790
rect 2176 -3858 2210 -3824
rect 2244 -3858 2278 -3824
rect 2312 -3858 2346 -3824
rect 2380 -3858 2414 -3824
rect 2448 -3858 2648 -3824
rect 2682 -3858 2716 -3824
rect 2750 -3858 2784 -3824
rect 2818 -3858 2852 -3824
rect 2886 -3858 2920 -3824
rect 2176 -3891 2920 -3858
rect 2176 -3892 2277 -3891
rect 2176 -3926 2210 -3892
rect 2244 -3926 2277 -3892
rect 2176 -3960 2277 -3926
rect 2819 -3892 2920 -3891
rect 2819 -3926 2852 -3892
rect 2886 -3926 2920 -3892
rect 2176 -3994 2210 -3960
rect 2244 -3994 2277 -3960
rect 2176 -4028 2277 -3994
rect 2176 -4062 2210 -4028
rect 2244 -4062 2277 -4028
rect 2176 -4262 2277 -4062
rect 2176 -4296 2210 -4262
rect 2244 -4296 2277 -4262
rect 2176 -4330 2277 -4296
rect 2176 -4364 2210 -4330
rect 2244 -4364 2277 -4330
rect 2176 -4398 2277 -4364
rect 2819 -3960 2920 -3926
rect 2819 -3994 2852 -3960
rect 2886 -3994 2920 -3960
rect 2819 -4028 2920 -3994
rect 2819 -4062 2852 -4028
rect 2886 -4062 2920 -4028
rect 2819 -4262 2920 -4062
rect 2819 -4296 2852 -4262
rect 2886 -4296 2920 -4262
rect 2819 -4330 2920 -4296
rect 2819 -4364 2852 -4330
rect 2886 -4364 2920 -4330
rect 2176 -4432 2210 -4398
rect 2244 -4432 2277 -4398
rect 2176 -4433 2277 -4432
rect 2819 -4398 2920 -4364
rect 2819 -4432 2852 -4398
rect 2886 -4432 2920 -4398
rect 2819 -4433 2920 -4432
rect 2176 -4466 2920 -4433
rect 2176 -4500 2210 -4466
rect 2244 -4500 2278 -4466
rect 2312 -4500 2346 -4466
rect 2380 -4500 2414 -4466
rect 2448 -4500 2648 -4466
rect 2682 -4500 2716 -4466
rect 2750 -4500 2784 -4466
rect 2818 -4500 2852 -4466
rect 2886 -4500 2920 -4466
rect 2176 -4534 2920 -4500
rect 2996 -3824 3740 -3790
rect 2996 -3858 3030 -3824
rect 3064 -3858 3098 -3824
rect 3132 -3858 3166 -3824
rect 3200 -3858 3234 -3824
rect 3268 -3858 3468 -3824
rect 3502 -3858 3536 -3824
rect 3570 -3858 3604 -3824
rect 3638 -3858 3672 -3824
rect 3706 -3858 3740 -3824
rect 2996 -3891 3740 -3858
rect 2996 -3892 3097 -3891
rect 2996 -3926 3030 -3892
rect 3064 -3926 3097 -3892
rect 2996 -3960 3097 -3926
rect 3639 -3892 3740 -3891
rect 3639 -3926 3672 -3892
rect 3706 -3926 3740 -3892
rect 2996 -3994 3030 -3960
rect 3064 -3994 3097 -3960
rect 2996 -4028 3097 -3994
rect 2996 -4062 3030 -4028
rect 3064 -4062 3097 -4028
rect 2996 -4262 3097 -4062
rect 2996 -4296 3030 -4262
rect 3064 -4296 3097 -4262
rect 2996 -4330 3097 -4296
rect 2996 -4364 3030 -4330
rect 3064 -4364 3097 -4330
rect 2996 -4398 3097 -4364
rect 3639 -3960 3740 -3926
rect 3639 -3994 3672 -3960
rect 3706 -3994 3740 -3960
rect 3639 -4028 3740 -3994
rect 3639 -4062 3672 -4028
rect 3706 -4062 3740 -4028
rect 3639 -4262 3740 -4062
rect 3639 -4296 3672 -4262
rect 3706 -4296 3740 -4262
rect 3639 -4330 3740 -4296
rect 3639 -4364 3672 -4330
rect 3706 -4364 3740 -4330
rect 2996 -4432 3030 -4398
rect 3064 -4432 3097 -4398
rect 2996 -4433 3097 -4432
rect 3639 -4398 3740 -4364
rect 3639 -4432 3672 -4398
rect 3706 -4432 3740 -4398
rect 3639 -4433 3740 -4432
rect 2996 -4466 3740 -4433
rect 2996 -4500 3030 -4466
rect 3064 -4500 3098 -4466
rect 3132 -4500 3166 -4466
rect 3200 -4500 3234 -4466
rect 3268 -4500 3468 -4466
rect 3502 -4500 3536 -4466
rect 3570 -4500 3604 -4466
rect 3638 -4500 3672 -4466
rect 3706 -4500 3740 -4466
rect 2996 -4534 3740 -4500
rect 3816 -3824 4560 -3790
rect 3816 -3858 3850 -3824
rect 3884 -3858 3918 -3824
rect 3952 -3858 3986 -3824
rect 4020 -3858 4054 -3824
rect 4088 -3858 4288 -3824
rect 4322 -3858 4356 -3824
rect 4390 -3858 4424 -3824
rect 4458 -3858 4492 -3824
rect 4526 -3858 4560 -3824
rect 3816 -3891 4560 -3858
rect 3816 -3892 3917 -3891
rect 3816 -3926 3850 -3892
rect 3884 -3926 3917 -3892
rect 3816 -3960 3917 -3926
rect 4459 -3892 4560 -3891
rect 4459 -3926 4492 -3892
rect 4526 -3926 4560 -3892
rect 3816 -3994 3850 -3960
rect 3884 -3994 3917 -3960
rect 3816 -4028 3917 -3994
rect 3816 -4062 3850 -4028
rect 3884 -4062 3917 -4028
rect 3816 -4262 3917 -4062
rect 3816 -4296 3850 -4262
rect 3884 -4296 3917 -4262
rect 3816 -4330 3917 -4296
rect 3816 -4364 3850 -4330
rect 3884 -4364 3917 -4330
rect 3816 -4398 3917 -4364
rect 4459 -3960 4560 -3926
rect 4459 -3994 4492 -3960
rect 4526 -3994 4560 -3960
rect 4459 -4028 4560 -3994
rect 4459 -4062 4492 -4028
rect 4526 -4062 4560 -4028
rect 4459 -4262 4560 -4062
rect 4459 -4296 4492 -4262
rect 4526 -4296 4560 -4262
rect 4459 -4330 4560 -4296
rect 4459 -4364 4492 -4330
rect 4526 -4364 4560 -4330
rect 3816 -4432 3850 -4398
rect 3884 -4432 3917 -4398
rect 3816 -4433 3917 -4432
rect 4459 -4398 4560 -4364
rect 4459 -4432 4492 -4398
rect 4526 -4432 4560 -4398
rect 4459 -4433 4560 -4432
rect 3816 -4466 4560 -4433
rect 3816 -4500 3850 -4466
rect 3884 -4500 3918 -4466
rect 3952 -4500 3986 -4466
rect 4020 -4500 4054 -4466
rect 4088 -4500 4288 -4466
rect 4322 -4500 4356 -4466
rect 4390 -4500 4424 -4466
rect 4458 -4500 4492 -4466
rect 4526 -4500 4560 -4466
rect 3816 -4534 4560 -4500
rect 4636 -3824 5380 -3790
rect 4636 -3858 4670 -3824
rect 4704 -3858 4738 -3824
rect 4772 -3858 4806 -3824
rect 4840 -3858 4874 -3824
rect 4908 -3858 5108 -3824
rect 5142 -3858 5176 -3824
rect 5210 -3858 5244 -3824
rect 5278 -3858 5312 -3824
rect 5346 -3858 5380 -3824
rect 4636 -3891 5380 -3858
rect 4636 -3892 4737 -3891
rect 4636 -3926 4670 -3892
rect 4704 -3926 4737 -3892
rect 4636 -3960 4737 -3926
rect 5279 -3892 5380 -3891
rect 5279 -3926 5312 -3892
rect 5346 -3926 5380 -3892
rect 4636 -3994 4670 -3960
rect 4704 -3994 4737 -3960
rect 4636 -4028 4737 -3994
rect 4636 -4062 4670 -4028
rect 4704 -4062 4737 -4028
rect 4636 -4262 4737 -4062
rect 4636 -4296 4670 -4262
rect 4704 -4296 4737 -4262
rect 4636 -4330 4737 -4296
rect 4636 -4364 4670 -4330
rect 4704 -4364 4737 -4330
rect 4636 -4398 4737 -4364
rect 5279 -3960 5380 -3926
rect 5279 -3994 5312 -3960
rect 5346 -3994 5380 -3960
rect 5279 -4028 5380 -3994
rect 5279 -4062 5312 -4028
rect 5346 -4062 5380 -4028
rect 5279 -4262 5380 -4062
rect 5279 -4296 5312 -4262
rect 5346 -4296 5380 -4262
rect 5279 -4330 5380 -4296
rect 5279 -4364 5312 -4330
rect 5346 -4364 5380 -4330
rect 4636 -4432 4670 -4398
rect 4704 -4432 4737 -4398
rect 4636 -4433 4737 -4432
rect 5279 -4398 5380 -4364
rect 5279 -4432 5312 -4398
rect 5346 -4432 5380 -4398
rect 5279 -4433 5380 -4432
rect 4636 -4466 5380 -4433
rect 4636 -4500 4670 -4466
rect 4704 -4500 4738 -4466
rect 4772 -4500 4806 -4466
rect 4840 -4500 4874 -4466
rect 4908 -4500 5108 -4466
rect 5142 -4500 5176 -4466
rect 5210 -4500 5244 -4466
rect 5278 -4500 5312 -4466
rect 5346 -4500 5380 -4466
rect 4636 -4534 5380 -4500
rect 5456 -3824 6200 -3790
rect 5456 -3858 5490 -3824
rect 5524 -3858 5558 -3824
rect 5592 -3858 5626 -3824
rect 5660 -3858 5694 -3824
rect 5728 -3858 5928 -3824
rect 5962 -3858 5996 -3824
rect 6030 -3858 6064 -3824
rect 6098 -3858 6132 -3824
rect 6166 -3858 6200 -3824
rect 5456 -3891 6200 -3858
rect 5456 -3892 5557 -3891
rect 5456 -3926 5490 -3892
rect 5524 -3926 5557 -3892
rect 5456 -3960 5557 -3926
rect 6099 -3892 6200 -3891
rect 6099 -3926 6132 -3892
rect 6166 -3926 6200 -3892
rect 5456 -3994 5490 -3960
rect 5524 -3994 5557 -3960
rect 5456 -4028 5557 -3994
rect 5456 -4062 5490 -4028
rect 5524 -4062 5557 -4028
rect 5456 -4262 5557 -4062
rect 5456 -4296 5490 -4262
rect 5524 -4296 5557 -4262
rect 5456 -4330 5557 -4296
rect 5456 -4364 5490 -4330
rect 5524 -4364 5557 -4330
rect 5456 -4398 5557 -4364
rect 6099 -3960 6200 -3926
rect 6099 -3994 6132 -3960
rect 6166 -3994 6200 -3960
rect 6099 -4028 6200 -3994
rect 6099 -4062 6132 -4028
rect 6166 -4062 6200 -4028
rect 6099 -4262 6200 -4062
rect 6099 -4296 6132 -4262
rect 6166 -4296 6200 -4262
rect 6099 -4330 6200 -4296
rect 6099 -4364 6132 -4330
rect 6166 -4364 6200 -4330
rect 5456 -4432 5490 -4398
rect 5524 -4432 5557 -4398
rect 5456 -4433 5557 -4432
rect 6099 -4398 6200 -4364
rect 6099 -4432 6132 -4398
rect 6166 -4432 6200 -4398
rect 6099 -4433 6200 -4432
rect 5456 -4466 6200 -4433
rect 5456 -4500 5490 -4466
rect 5524 -4500 5558 -4466
rect 5592 -4500 5626 -4466
rect 5660 -4500 5694 -4466
rect 5728 -4500 5928 -4466
rect 5962 -4500 5996 -4466
rect 6030 -4500 6064 -4466
rect 6098 -4500 6132 -4466
rect 6166 -4500 6200 -4466
rect 5456 -4534 6200 -4500
rect 6276 -3824 7020 -3790
rect 6276 -3858 6310 -3824
rect 6344 -3858 6378 -3824
rect 6412 -3858 6446 -3824
rect 6480 -3858 6514 -3824
rect 6548 -3858 6748 -3824
rect 6782 -3858 6816 -3824
rect 6850 -3858 6884 -3824
rect 6918 -3858 6952 -3824
rect 6986 -3858 7020 -3824
rect 6276 -3891 7020 -3858
rect 6276 -3892 6377 -3891
rect 6276 -3926 6310 -3892
rect 6344 -3926 6377 -3892
rect 6276 -3960 6377 -3926
rect 6919 -3892 7020 -3891
rect 6919 -3926 6952 -3892
rect 6986 -3926 7020 -3892
rect 6276 -3994 6310 -3960
rect 6344 -3994 6377 -3960
rect 6276 -4028 6377 -3994
rect 6276 -4062 6310 -4028
rect 6344 -4062 6377 -4028
rect 6276 -4262 6377 -4062
rect 6276 -4296 6310 -4262
rect 6344 -4296 6377 -4262
rect 6276 -4330 6377 -4296
rect 6276 -4364 6310 -4330
rect 6344 -4364 6377 -4330
rect 6276 -4398 6377 -4364
rect 6919 -3960 7020 -3926
rect 6919 -3994 6952 -3960
rect 6986 -3994 7020 -3960
rect 6919 -4028 7020 -3994
rect 6919 -4062 6952 -4028
rect 6986 -4062 7020 -4028
rect 6919 -4262 7020 -4062
rect 6919 -4296 6952 -4262
rect 6986 -4296 7020 -4262
rect 6919 -4330 7020 -4296
rect 6919 -4364 6952 -4330
rect 6986 -4364 7020 -4330
rect 6276 -4432 6310 -4398
rect 6344 -4432 6377 -4398
rect 6276 -4433 6377 -4432
rect 6919 -4398 7020 -4364
rect 6919 -4432 6952 -4398
rect 6986 -4432 7020 -4398
rect 6919 -4433 7020 -4432
rect 6276 -4466 7020 -4433
rect 6276 -4500 6310 -4466
rect 6344 -4500 6378 -4466
rect 6412 -4500 6446 -4466
rect 6480 -4500 6514 -4466
rect 6548 -4500 6748 -4466
rect 6782 -4500 6816 -4466
rect 6850 -4500 6884 -4466
rect 6918 -4500 6952 -4466
rect 6986 -4500 7020 -4466
rect 6276 -4534 7020 -4500
<< nsubdiff >>
rect 7630 6240 7730 6270
rect 7630 4300 7660 6240
rect 7700 4300 7730 6240
rect 7630 4270 7730 4300
rect 7630 4030 7730 4060
rect 7630 2090 7660 4030
rect 7700 2090 7730 4030
rect 7630 2060 7730 2090
rect -941 -697 -523 -673
rect -941 -731 -917 -697
rect -883 -731 -849 -697
rect -815 -731 -649 -697
rect -615 -731 -581 -697
rect -547 -731 -523 -697
rect -941 -745 -523 -731
rect -941 -765 -869 -745
rect -941 -799 -917 -765
rect -883 -799 -869 -765
rect -941 -965 -869 -799
rect -595 -765 -523 -745
rect -595 -799 -581 -765
rect -547 -799 -523 -765
rect -941 -999 -917 -965
rect -883 -999 -869 -965
rect -941 -1019 -869 -999
rect -595 -965 -523 -799
rect -595 -999 -581 -965
rect -547 -999 -523 -965
rect -595 -1019 -523 -999
rect -941 -1033 -523 -1019
rect -941 -1067 -917 -1033
rect -883 -1067 -849 -1033
rect -815 -1067 -649 -1033
rect -615 -1067 -581 -1033
rect -547 -1067 -523 -1033
rect -941 -1091 -523 -1067
rect -121 -697 297 -673
rect -121 -731 -97 -697
rect -63 -731 -29 -697
rect 5 -731 171 -697
rect 205 -731 239 -697
rect 273 -731 297 -697
rect -121 -745 297 -731
rect -121 -765 -49 -745
rect -121 -799 -97 -765
rect -63 -799 -49 -765
rect -121 -965 -49 -799
rect 225 -765 297 -745
rect 225 -799 239 -765
rect 273 -799 297 -765
rect -121 -999 -97 -965
rect -63 -999 -49 -965
rect -121 -1019 -49 -999
rect 225 -965 297 -799
rect 225 -999 239 -965
rect 273 -999 297 -965
rect 225 -1019 297 -999
rect -121 -1033 297 -1019
rect -121 -1067 -97 -1033
rect -63 -1067 -29 -1033
rect 5 -1067 171 -1033
rect 205 -1067 239 -1033
rect 273 -1067 297 -1033
rect -121 -1091 297 -1067
rect 699 -697 1117 -673
rect 699 -731 723 -697
rect 757 -731 791 -697
rect 825 -731 991 -697
rect 1025 -731 1059 -697
rect 1093 -731 1117 -697
rect 699 -745 1117 -731
rect 699 -765 771 -745
rect 699 -799 723 -765
rect 757 -799 771 -765
rect 699 -965 771 -799
rect 1045 -765 1117 -745
rect 1045 -799 1059 -765
rect 1093 -799 1117 -765
rect 699 -999 723 -965
rect 757 -999 771 -965
rect 699 -1019 771 -999
rect 1045 -965 1117 -799
rect 1045 -999 1059 -965
rect 1093 -999 1117 -965
rect 1045 -1019 1117 -999
rect 699 -1033 1117 -1019
rect 699 -1067 723 -1033
rect 757 -1067 791 -1033
rect 825 -1067 991 -1033
rect 1025 -1067 1059 -1033
rect 1093 -1067 1117 -1033
rect 699 -1091 1117 -1067
rect 1519 -697 1937 -673
rect 1519 -731 1543 -697
rect 1577 -731 1611 -697
rect 1645 -731 1811 -697
rect 1845 -731 1879 -697
rect 1913 -731 1937 -697
rect 1519 -745 1937 -731
rect 1519 -765 1591 -745
rect 1519 -799 1543 -765
rect 1577 -799 1591 -765
rect 1519 -965 1591 -799
rect 1865 -765 1937 -745
rect 1865 -799 1879 -765
rect 1913 -799 1937 -765
rect 1519 -999 1543 -965
rect 1577 -999 1591 -965
rect 1519 -1019 1591 -999
rect 1865 -965 1937 -799
rect 1865 -999 1879 -965
rect 1913 -999 1937 -965
rect 1865 -1019 1937 -999
rect 1519 -1033 1937 -1019
rect 1519 -1067 1543 -1033
rect 1577 -1067 1611 -1033
rect 1645 -1067 1811 -1033
rect 1845 -1067 1879 -1033
rect 1913 -1067 1937 -1033
rect 1519 -1091 1937 -1067
rect 2339 -697 2757 -673
rect 2339 -731 2363 -697
rect 2397 -731 2431 -697
rect 2465 -731 2631 -697
rect 2665 -731 2699 -697
rect 2733 -731 2757 -697
rect 2339 -745 2757 -731
rect 2339 -765 2411 -745
rect 2339 -799 2363 -765
rect 2397 -799 2411 -765
rect 2339 -965 2411 -799
rect 2685 -765 2757 -745
rect 2685 -799 2699 -765
rect 2733 -799 2757 -765
rect 2339 -999 2363 -965
rect 2397 -999 2411 -965
rect 2339 -1019 2411 -999
rect 2685 -965 2757 -799
rect 2685 -999 2699 -965
rect 2733 -999 2757 -965
rect 2685 -1019 2757 -999
rect 2339 -1033 2757 -1019
rect 2339 -1067 2363 -1033
rect 2397 -1067 2431 -1033
rect 2465 -1067 2631 -1033
rect 2665 -1067 2699 -1033
rect 2733 -1067 2757 -1033
rect 2339 -1091 2757 -1067
rect 3159 -697 3577 -673
rect 3159 -731 3183 -697
rect 3217 -731 3251 -697
rect 3285 -731 3451 -697
rect 3485 -731 3519 -697
rect 3553 -731 3577 -697
rect 3159 -745 3577 -731
rect 3159 -765 3231 -745
rect 3159 -799 3183 -765
rect 3217 -799 3231 -765
rect 3159 -965 3231 -799
rect 3505 -765 3577 -745
rect 3505 -799 3519 -765
rect 3553 -799 3577 -765
rect 3159 -999 3183 -965
rect 3217 -999 3231 -965
rect 3159 -1019 3231 -999
rect 3505 -965 3577 -799
rect 3505 -999 3519 -965
rect 3553 -999 3577 -965
rect 3505 -1019 3577 -999
rect 3159 -1033 3577 -1019
rect 3159 -1067 3183 -1033
rect 3217 -1067 3251 -1033
rect 3285 -1067 3451 -1033
rect 3485 -1067 3519 -1033
rect 3553 -1067 3577 -1033
rect 3159 -1091 3577 -1067
rect 3979 -697 4397 -673
rect 3979 -731 4003 -697
rect 4037 -731 4071 -697
rect 4105 -731 4271 -697
rect 4305 -731 4339 -697
rect 4373 -731 4397 -697
rect 3979 -745 4397 -731
rect 3979 -765 4051 -745
rect 3979 -799 4003 -765
rect 4037 -799 4051 -765
rect 3979 -965 4051 -799
rect 4325 -765 4397 -745
rect 4325 -799 4339 -765
rect 4373 -799 4397 -765
rect 3979 -999 4003 -965
rect 4037 -999 4051 -965
rect 3979 -1019 4051 -999
rect 4325 -965 4397 -799
rect 4325 -999 4339 -965
rect 4373 -999 4397 -965
rect 4325 -1019 4397 -999
rect 3979 -1033 4397 -1019
rect 3979 -1067 4003 -1033
rect 4037 -1067 4071 -1033
rect 4105 -1067 4271 -1033
rect 4305 -1067 4339 -1033
rect 4373 -1067 4397 -1033
rect 3979 -1091 4397 -1067
rect 4799 -697 5217 -673
rect 4799 -731 4823 -697
rect 4857 -731 4891 -697
rect 4925 -731 5091 -697
rect 5125 -731 5159 -697
rect 5193 -731 5217 -697
rect 4799 -745 5217 -731
rect 4799 -765 4871 -745
rect 4799 -799 4823 -765
rect 4857 -799 4871 -765
rect 4799 -965 4871 -799
rect 5145 -765 5217 -745
rect 5145 -799 5159 -765
rect 5193 -799 5217 -765
rect 4799 -999 4823 -965
rect 4857 -999 4871 -965
rect 4799 -1019 4871 -999
rect 5145 -965 5217 -799
rect 5145 -999 5159 -965
rect 5193 -999 5217 -965
rect 5145 -1019 5217 -999
rect 4799 -1033 5217 -1019
rect 4799 -1067 4823 -1033
rect 4857 -1067 4891 -1033
rect 4925 -1067 5091 -1033
rect 5125 -1067 5159 -1033
rect 5193 -1067 5217 -1033
rect 4799 -1091 5217 -1067
rect 5619 -697 6037 -673
rect 5619 -731 5643 -697
rect 5677 -731 5711 -697
rect 5745 -731 5911 -697
rect 5945 -731 5979 -697
rect 6013 -731 6037 -697
rect 5619 -745 6037 -731
rect 5619 -765 5691 -745
rect 5619 -799 5643 -765
rect 5677 -799 5691 -765
rect 5619 -965 5691 -799
rect 5965 -765 6037 -745
rect 5965 -799 5979 -765
rect 6013 -799 6037 -765
rect 5619 -999 5643 -965
rect 5677 -999 5691 -965
rect 5619 -1019 5691 -999
rect 5965 -965 6037 -799
rect 5965 -999 5979 -965
rect 6013 -999 6037 -965
rect 5965 -1019 6037 -999
rect 5619 -1033 6037 -1019
rect 5619 -1067 5643 -1033
rect 5677 -1067 5711 -1033
rect 5745 -1067 5911 -1033
rect 5945 -1067 5979 -1033
rect 6013 -1067 6037 -1033
rect 5619 -1091 6037 -1067
rect 6439 -697 6857 -673
rect 6439 -731 6463 -697
rect 6497 -731 6531 -697
rect 6565 -731 6731 -697
rect 6765 -731 6799 -697
rect 6833 -731 6857 -697
rect 6439 -745 6857 -731
rect 6439 -765 6511 -745
rect 6439 -799 6463 -765
rect 6497 -799 6511 -765
rect 6439 -965 6511 -799
rect 6785 -765 6857 -745
rect 6785 -799 6799 -765
rect 6833 -799 6857 -765
rect 6439 -999 6463 -965
rect 6497 -999 6511 -965
rect 6439 -1019 6511 -999
rect 6785 -965 6857 -799
rect 6785 -999 6799 -965
rect 6833 -999 6857 -965
rect 6785 -1019 6857 -999
rect 6439 -1033 6857 -1019
rect 6439 -1067 6463 -1033
rect 6497 -1067 6531 -1033
rect 6565 -1067 6731 -1033
rect 6765 -1067 6799 -1033
rect 6833 -1067 6857 -1033
rect 6439 -1091 6857 -1067
rect 7289 -697 7707 -673
rect 7289 -731 7313 -697
rect 7347 -731 7381 -697
rect 7415 -731 7581 -697
rect 7615 -731 7649 -697
rect 7683 -731 7707 -697
rect 7289 -745 7707 -731
rect 7289 -765 7361 -745
rect 7289 -799 7313 -765
rect 7347 -799 7361 -765
rect 7289 -965 7361 -799
rect 7635 -765 7707 -745
rect 7635 -799 7649 -765
rect 7683 -799 7707 -765
rect 7289 -999 7313 -965
rect 7347 -999 7361 -965
rect 7289 -1019 7361 -999
rect 7635 -965 7707 -799
rect 7635 -999 7649 -965
rect 7683 -999 7707 -965
rect 7635 -1019 7707 -999
rect 7289 -1033 7707 -1019
rect 7289 -1067 7313 -1033
rect 7347 -1067 7381 -1033
rect 7415 -1067 7581 -1033
rect 7615 -1067 7649 -1033
rect 7683 -1067 7707 -1033
rect 7289 -1091 7707 -1067
rect -941 -1517 -523 -1493
rect -941 -1551 -917 -1517
rect -883 -1551 -849 -1517
rect -815 -1551 -649 -1517
rect -615 -1551 -581 -1517
rect -547 -1551 -523 -1517
rect -941 -1565 -523 -1551
rect -941 -1585 -869 -1565
rect -941 -1619 -917 -1585
rect -883 -1619 -869 -1585
rect -941 -1785 -869 -1619
rect -595 -1585 -523 -1565
rect -595 -1619 -581 -1585
rect -547 -1619 -523 -1585
rect -941 -1819 -917 -1785
rect -883 -1819 -869 -1785
rect -941 -1839 -869 -1819
rect -595 -1785 -523 -1619
rect -595 -1819 -581 -1785
rect -547 -1819 -523 -1785
rect -595 -1839 -523 -1819
rect -941 -1853 -523 -1839
rect -941 -1887 -917 -1853
rect -883 -1887 -849 -1853
rect -815 -1887 -649 -1853
rect -615 -1887 -581 -1853
rect -547 -1887 -523 -1853
rect -941 -1911 -523 -1887
rect -121 -1517 297 -1493
rect -121 -1551 -97 -1517
rect -63 -1551 -29 -1517
rect 5 -1551 171 -1517
rect 205 -1551 239 -1517
rect 273 -1551 297 -1517
rect -121 -1565 297 -1551
rect -121 -1585 -49 -1565
rect -121 -1619 -97 -1585
rect -63 -1619 -49 -1585
rect -121 -1785 -49 -1619
rect 225 -1585 297 -1565
rect 225 -1619 239 -1585
rect 273 -1619 297 -1585
rect -121 -1819 -97 -1785
rect -63 -1819 -49 -1785
rect -121 -1839 -49 -1819
rect 225 -1785 297 -1619
rect 225 -1819 239 -1785
rect 273 -1819 297 -1785
rect 225 -1839 297 -1819
rect -121 -1853 297 -1839
rect -121 -1887 -97 -1853
rect -63 -1887 -29 -1853
rect 5 -1887 171 -1853
rect 205 -1887 239 -1853
rect 273 -1887 297 -1853
rect -121 -1911 297 -1887
rect 699 -1517 1117 -1493
rect 699 -1551 723 -1517
rect 757 -1551 791 -1517
rect 825 -1551 991 -1517
rect 1025 -1551 1059 -1517
rect 1093 -1551 1117 -1517
rect 699 -1565 1117 -1551
rect 699 -1585 771 -1565
rect 699 -1619 723 -1585
rect 757 -1619 771 -1585
rect 699 -1785 771 -1619
rect 1045 -1585 1117 -1565
rect 1045 -1619 1059 -1585
rect 1093 -1619 1117 -1585
rect 699 -1819 723 -1785
rect 757 -1819 771 -1785
rect 699 -1839 771 -1819
rect 1045 -1785 1117 -1619
rect 1045 -1819 1059 -1785
rect 1093 -1819 1117 -1785
rect 1045 -1839 1117 -1819
rect 699 -1853 1117 -1839
rect 699 -1887 723 -1853
rect 757 -1887 791 -1853
rect 825 -1887 991 -1853
rect 1025 -1887 1059 -1853
rect 1093 -1887 1117 -1853
rect 699 -1911 1117 -1887
rect 1519 -1517 1937 -1493
rect 1519 -1551 1543 -1517
rect 1577 -1551 1611 -1517
rect 1645 -1551 1811 -1517
rect 1845 -1551 1879 -1517
rect 1913 -1551 1937 -1517
rect 1519 -1565 1937 -1551
rect 1519 -1585 1591 -1565
rect 1519 -1619 1543 -1585
rect 1577 -1619 1591 -1585
rect 1519 -1785 1591 -1619
rect 1865 -1585 1937 -1565
rect 1865 -1619 1879 -1585
rect 1913 -1619 1937 -1585
rect 1519 -1819 1543 -1785
rect 1577 -1819 1591 -1785
rect 1519 -1839 1591 -1819
rect 1865 -1785 1937 -1619
rect 1865 -1819 1879 -1785
rect 1913 -1819 1937 -1785
rect 1865 -1839 1937 -1819
rect 1519 -1853 1937 -1839
rect 1519 -1887 1543 -1853
rect 1577 -1887 1611 -1853
rect 1645 -1887 1811 -1853
rect 1845 -1887 1879 -1853
rect 1913 -1887 1937 -1853
rect 1519 -1911 1937 -1887
rect 2339 -1517 2757 -1493
rect 2339 -1551 2363 -1517
rect 2397 -1551 2431 -1517
rect 2465 -1551 2631 -1517
rect 2665 -1551 2699 -1517
rect 2733 -1551 2757 -1517
rect 2339 -1565 2757 -1551
rect 2339 -1585 2411 -1565
rect 2339 -1619 2363 -1585
rect 2397 -1619 2411 -1585
rect 2339 -1785 2411 -1619
rect 2685 -1585 2757 -1565
rect 2685 -1619 2699 -1585
rect 2733 -1619 2757 -1585
rect 2339 -1819 2363 -1785
rect 2397 -1819 2411 -1785
rect 2339 -1839 2411 -1819
rect 2685 -1785 2757 -1619
rect 2685 -1819 2699 -1785
rect 2733 -1819 2757 -1785
rect 2685 -1839 2757 -1819
rect 2339 -1853 2757 -1839
rect 2339 -1887 2363 -1853
rect 2397 -1887 2431 -1853
rect 2465 -1887 2631 -1853
rect 2665 -1887 2699 -1853
rect 2733 -1887 2757 -1853
rect 2339 -1911 2757 -1887
rect 3159 -1517 3577 -1493
rect 3159 -1551 3183 -1517
rect 3217 -1551 3251 -1517
rect 3285 -1551 3451 -1517
rect 3485 -1551 3519 -1517
rect 3553 -1551 3577 -1517
rect 3159 -1565 3577 -1551
rect 3159 -1585 3231 -1565
rect 3159 -1619 3183 -1585
rect 3217 -1619 3231 -1585
rect 3159 -1785 3231 -1619
rect 3505 -1585 3577 -1565
rect 3505 -1619 3519 -1585
rect 3553 -1619 3577 -1585
rect 3159 -1819 3183 -1785
rect 3217 -1819 3231 -1785
rect 3159 -1839 3231 -1819
rect 3505 -1785 3577 -1619
rect 3505 -1819 3519 -1785
rect 3553 -1819 3577 -1785
rect 3505 -1839 3577 -1819
rect 3159 -1853 3577 -1839
rect 3159 -1887 3183 -1853
rect 3217 -1887 3251 -1853
rect 3285 -1887 3451 -1853
rect 3485 -1887 3519 -1853
rect 3553 -1887 3577 -1853
rect 3159 -1911 3577 -1887
rect 3979 -1517 4397 -1493
rect 3979 -1551 4003 -1517
rect 4037 -1551 4071 -1517
rect 4105 -1551 4271 -1517
rect 4305 -1551 4339 -1517
rect 4373 -1551 4397 -1517
rect 3979 -1565 4397 -1551
rect 3979 -1585 4051 -1565
rect 3979 -1619 4003 -1585
rect 4037 -1619 4051 -1585
rect 3979 -1785 4051 -1619
rect 4325 -1585 4397 -1565
rect 4325 -1619 4339 -1585
rect 4373 -1619 4397 -1585
rect 3979 -1819 4003 -1785
rect 4037 -1819 4051 -1785
rect 3979 -1839 4051 -1819
rect 4325 -1785 4397 -1619
rect 4325 -1819 4339 -1785
rect 4373 -1819 4397 -1785
rect 4325 -1839 4397 -1819
rect 3979 -1853 4397 -1839
rect 3979 -1887 4003 -1853
rect 4037 -1887 4071 -1853
rect 4105 -1887 4271 -1853
rect 4305 -1887 4339 -1853
rect 4373 -1887 4397 -1853
rect 3979 -1911 4397 -1887
rect 4799 -1517 5217 -1493
rect 4799 -1551 4823 -1517
rect 4857 -1551 4891 -1517
rect 4925 -1551 5091 -1517
rect 5125 -1551 5159 -1517
rect 5193 -1551 5217 -1517
rect 4799 -1565 5217 -1551
rect 4799 -1585 4871 -1565
rect 4799 -1619 4823 -1585
rect 4857 -1619 4871 -1585
rect 4799 -1785 4871 -1619
rect 5145 -1585 5217 -1565
rect 5145 -1619 5159 -1585
rect 5193 -1619 5217 -1585
rect 4799 -1819 4823 -1785
rect 4857 -1819 4871 -1785
rect 4799 -1839 4871 -1819
rect 5145 -1785 5217 -1619
rect 5145 -1819 5159 -1785
rect 5193 -1819 5217 -1785
rect 5145 -1839 5217 -1819
rect 4799 -1853 5217 -1839
rect 4799 -1887 4823 -1853
rect 4857 -1887 4891 -1853
rect 4925 -1887 5091 -1853
rect 5125 -1887 5159 -1853
rect 5193 -1887 5217 -1853
rect 4799 -1911 5217 -1887
rect 5619 -1517 6037 -1493
rect 5619 -1551 5643 -1517
rect 5677 -1551 5711 -1517
rect 5745 -1551 5911 -1517
rect 5945 -1551 5979 -1517
rect 6013 -1551 6037 -1517
rect 5619 -1565 6037 -1551
rect 5619 -1585 5691 -1565
rect 5619 -1619 5643 -1585
rect 5677 -1619 5691 -1585
rect 5619 -1785 5691 -1619
rect 5965 -1585 6037 -1565
rect 5965 -1619 5979 -1585
rect 6013 -1619 6037 -1585
rect 5619 -1819 5643 -1785
rect 5677 -1819 5691 -1785
rect 5619 -1839 5691 -1819
rect 5965 -1785 6037 -1619
rect 5965 -1819 5979 -1785
rect 6013 -1819 6037 -1785
rect 5965 -1839 6037 -1819
rect 5619 -1853 6037 -1839
rect 5619 -1887 5643 -1853
rect 5677 -1887 5711 -1853
rect 5745 -1887 5911 -1853
rect 5945 -1887 5979 -1853
rect 6013 -1887 6037 -1853
rect 5619 -1911 6037 -1887
rect 6439 -1517 6857 -1493
rect 6439 -1551 6463 -1517
rect 6497 -1551 6531 -1517
rect 6565 -1551 6731 -1517
rect 6765 -1551 6799 -1517
rect 6833 -1551 6857 -1517
rect 6439 -1565 6857 -1551
rect 6439 -1585 6511 -1565
rect 6439 -1619 6463 -1585
rect 6497 -1619 6511 -1585
rect 6439 -1785 6511 -1619
rect 6785 -1585 6857 -1565
rect 6785 -1619 6799 -1585
rect 6833 -1619 6857 -1585
rect 6439 -1819 6463 -1785
rect 6497 -1819 6511 -1785
rect 6439 -1839 6511 -1819
rect 6785 -1785 6857 -1619
rect 6785 -1819 6799 -1785
rect 6833 -1819 6857 -1785
rect 6785 -1839 6857 -1819
rect 6439 -1853 6857 -1839
rect 6439 -1887 6463 -1853
rect 6497 -1887 6531 -1853
rect 6565 -1887 6731 -1853
rect 6765 -1887 6799 -1853
rect 6833 -1887 6857 -1853
rect 6439 -1911 6857 -1887
rect -941 -2337 -523 -2313
rect -941 -2371 -917 -2337
rect -883 -2371 -849 -2337
rect -815 -2371 -649 -2337
rect -615 -2371 -581 -2337
rect -547 -2371 -523 -2337
rect -941 -2385 -523 -2371
rect -941 -2405 -869 -2385
rect -941 -2439 -917 -2405
rect -883 -2439 -869 -2405
rect -941 -2605 -869 -2439
rect -595 -2405 -523 -2385
rect -595 -2439 -581 -2405
rect -547 -2439 -523 -2405
rect -941 -2639 -917 -2605
rect -883 -2639 -869 -2605
rect -941 -2659 -869 -2639
rect -595 -2605 -523 -2439
rect -595 -2639 -581 -2605
rect -547 -2639 -523 -2605
rect -595 -2659 -523 -2639
rect -941 -2673 -523 -2659
rect -941 -2707 -917 -2673
rect -883 -2707 -849 -2673
rect -815 -2707 -649 -2673
rect -615 -2707 -581 -2673
rect -547 -2707 -523 -2673
rect -941 -2731 -523 -2707
rect -121 -2337 297 -2313
rect -121 -2371 -97 -2337
rect -63 -2371 -29 -2337
rect 5 -2371 171 -2337
rect 205 -2371 239 -2337
rect 273 -2371 297 -2337
rect -121 -2385 297 -2371
rect -121 -2405 -49 -2385
rect -121 -2439 -97 -2405
rect -63 -2439 -49 -2405
rect -121 -2605 -49 -2439
rect 225 -2405 297 -2385
rect 225 -2439 239 -2405
rect 273 -2439 297 -2405
rect -121 -2639 -97 -2605
rect -63 -2639 -49 -2605
rect -121 -2659 -49 -2639
rect 225 -2605 297 -2439
rect 225 -2639 239 -2605
rect 273 -2639 297 -2605
rect 225 -2659 297 -2639
rect -121 -2673 297 -2659
rect -121 -2707 -97 -2673
rect -63 -2707 -29 -2673
rect 5 -2707 171 -2673
rect 205 -2707 239 -2673
rect 273 -2707 297 -2673
rect -121 -2731 297 -2707
rect 699 -2337 1117 -2313
rect 699 -2371 723 -2337
rect 757 -2371 791 -2337
rect 825 -2371 991 -2337
rect 1025 -2371 1059 -2337
rect 1093 -2371 1117 -2337
rect 699 -2385 1117 -2371
rect 699 -2405 771 -2385
rect 699 -2439 723 -2405
rect 757 -2439 771 -2405
rect 699 -2605 771 -2439
rect 1045 -2405 1117 -2385
rect 1045 -2439 1059 -2405
rect 1093 -2439 1117 -2405
rect 699 -2639 723 -2605
rect 757 -2639 771 -2605
rect 699 -2659 771 -2639
rect 1045 -2605 1117 -2439
rect 1045 -2639 1059 -2605
rect 1093 -2639 1117 -2605
rect 1045 -2659 1117 -2639
rect 699 -2673 1117 -2659
rect 699 -2707 723 -2673
rect 757 -2707 791 -2673
rect 825 -2707 991 -2673
rect 1025 -2707 1059 -2673
rect 1093 -2707 1117 -2673
rect 699 -2731 1117 -2707
rect 1519 -2337 1937 -2313
rect 1519 -2371 1543 -2337
rect 1577 -2371 1611 -2337
rect 1645 -2371 1811 -2337
rect 1845 -2371 1879 -2337
rect 1913 -2371 1937 -2337
rect 1519 -2385 1937 -2371
rect 1519 -2405 1591 -2385
rect 1519 -2439 1543 -2405
rect 1577 -2439 1591 -2405
rect 1519 -2605 1591 -2439
rect 1865 -2405 1937 -2385
rect 1865 -2439 1879 -2405
rect 1913 -2439 1937 -2405
rect 1519 -2639 1543 -2605
rect 1577 -2639 1591 -2605
rect 1519 -2659 1591 -2639
rect 1865 -2605 1937 -2439
rect 1865 -2639 1879 -2605
rect 1913 -2639 1937 -2605
rect 1865 -2659 1937 -2639
rect 1519 -2673 1937 -2659
rect 1519 -2707 1543 -2673
rect 1577 -2707 1611 -2673
rect 1645 -2707 1811 -2673
rect 1845 -2707 1879 -2673
rect 1913 -2707 1937 -2673
rect 1519 -2731 1937 -2707
rect 2339 -2337 2757 -2313
rect 2339 -2371 2363 -2337
rect 2397 -2371 2431 -2337
rect 2465 -2371 2631 -2337
rect 2665 -2371 2699 -2337
rect 2733 -2371 2757 -2337
rect 2339 -2385 2757 -2371
rect 2339 -2405 2411 -2385
rect 2339 -2439 2363 -2405
rect 2397 -2439 2411 -2405
rect 2339 -2605 2411 -2439
rect 2685 -2405 2757 -2385
rect 2685 -2439 2699 -2405
rect 2733 -2439 2757 -2405
rect 2339 -2639 2363 -2605
rect 2397 -2639 2411 -2605
rect 2339 -2659 2411 -2639
rect 2685 -2605 2757 -2439
rect 2685 -2639 2699 -2605
rect 2733 -2639 2757 -2605
rect 2685 -2659 2757 -2639
rect 2339 -2673 2757 -2659
rect 2339 -2707 2363 -2673
rect 2397 -2707 2431 -2673
rect 2465 -2707 2631 -2673
rect 2665 -2707 2699 -2673
rect 2733 -2707 2757 -2673
rect 2339 -2731 2757 -2707
rect 3159 -2337 3577 -2313
rect 3159 -2371 3183 -2337
rect 3217 -2371 3251 -2337
rect 3285 -2371 3451 -2337
rect 3485 -2371 3519 -2337
rect 3553 -2371 3577 -2337
rect 3159 -2385 3577 -2371
rect 3159 -2405 3231 -2385
rect 3159 -2439 3183 -2405
rect 3217 -2439 3231 -2405
rect 3159 -2605 3231 -2439
rect 3505 -2405 3577 -2385
rect 3505 -2439 3519 -2405
rect 3553 -2439 3577 -2405
rect 3159 -2639 3183 -2605
rect 3217 -2639 3231 -2605
rect 3159 -2659 3231 -2639
rect 3505 -2605 3577 -2439
rect 3505 -2639 3519 -2605
rect 3553 -2639 3577 -2605
rect 3505 -2659 3577 -2639
rect 3159 -2673 3577 -2659
rect 3159 -2707 3183 -2673
rect 3217 -2707 3251 -2673
rect 3285 -2707 3451 -2673
rect 3485 -2707 3519 -2673
rect 3553 -2707 3577 -2673
rect 3159 -2731 3577 -2707
rect 3979 -2337 4397 -2313
rect 3979 -2371 4003 -2337
rect 4037 -2371 4071 -2337
rect 4105 -2371 4271 -2337
rect 4305 -2371 4339 -2337
rect 4373 -2371 4397 -2337
rect 3979 -2385 4397 -2371
rect 3979 -2405 4051 -2385
rect 3979 -2439 4003 -2405
rect 4037 -2439 4051 -2405
rect 3979 -2605 4051 -2439
rect 4325 -2405 4397 -2385
rect 4325 -2439 4339 -2405
rect 4373 -2439 4397 -2405
rect 3979 -2639 4003 -2605
rect 4037 -2639 4051 -2605
rect 3979 -2659 4051 -2639
rect 4325 -2605 4397 -2439
rect 4325 -2639 4339 -2605
rect 4373 -2639 4397 -2605
rect 4325 -2659 4397 -2639
rect 3979 -2673 4397 -2659
rect 3979 -2707 4003 -2673
rect 4037 -2707 4071 -2673
rect 4105 -2707 4271 -2673
rect 4305 -2707 4339 -2673
rect 4373 -2707 4397 -2673
rect 3979 -2731 4397 -2707
rect 4799 -2337 5217 -2313
rect 4799 -2371 4823 -2337
rect 4857 -2371 4891 -2337
rect 4925 -2371 5091 -2337
rect 5125 -2371 5159 -2337
rect 5193 -2371 5217 -2337
rect 4799 -2385 5217 -2371
rect 4799 -2405 4871 -2385
rect 4799 -2439 4823 -2405
rect 4857 -2439 4871 -2405
rect 4799 -2605 4871 -2439
rect 5145 -2405 5217 -2385
rect 5145 -2439 5159 -2405
rect 5193 -2439 5217 -2405
rect 4799 -2639 4823 -2605
rect 4857 -2639 4871 -2605
rect 4799 -2659 4871 -2639
rect 5145 -2605 5217 -2439
rect 5145 -2639 5159 -2605
rect 5193 -2639 5217 -2605
rect 5145 -2659 5217 -2639
rect 4799 -2673 5217 -2659
rect 4799 -2707 4823 -2673
rect 4857 -2707 4891 -2673
rect 4925 -2707 5091 -2673
rect 5125 -2707 5159 -2673
rect 5193 -2707 5217 -2673
rect 4799 -2731 5217 -2707
rect 5619 -2337 6037 -2313
rect 5619 -2371 5643 -2337
rect 5677 -2371 5711 -2337
rect 5745 -2371 5911 -2337
rect 5945 -2371 5979 -2337
rect 6013 -2371 6037 -2337
rect 5619 -2385 6037 -2371
rect 5619 -2405 5691 -2385
rect 5619 -2439 5643 -2405
rect 5677 -2439 5691 -2405
rect 5619 -2605 5691 -2439
rect 5965 -2405 6037 -2385
rect 5965 -2439 5979 -2405
rect 6013 -2439 6037 -2405
rect 5619 -2639 5643 -2605
rect 5677 -2639 5691 -2605
rect 5619 -2659 5691 -2639
rect 5965 -2605 6037 -2439
rect 5965 -2639 5979 -2605
rect 6013 -2639 6037 -2605
rect 5965 -2659 6037 -2639
rect 5619 -2673 6037 -2659
rect 5619 -2707 5643 -2673
rect 5677 -2707 5711 -2673
rect 5745 -2707 5911 -2673
rect 5945 -2707 5979 -2673
rect 6013 -2707 6037 -2673
rect 5619 -2731 6037 -2707
rect 6439 -2337 6857 -2313
rect 6439 -2371 6463 -2337
rect 6497 -2371 6531 -2337
rect 6565 -2371 6731 -2337
rect 6765 -2371 6799 -2337
rect 6833 -2371 6857 -2337
rect 6439 -2385 6857 -2371
rect 6439 -2405 6511 -2385
rect 6439 -2439 6463 -2405
rect 6497 -2439 6511 -2405
rect 6439 -2605 6511 -2439
rect 6785 -2405 6857 -2385
rect 6785 -2439 6799 -2405
rect 6833 -2439 6857 -2405
rect 6439 -2639 6463 -2605
rect 6497 -2639 6511 -2605
rect 6439 -2659 6511 -2639
rect 6785 -2605 6857 -2439
rect 6785 -2639 6799 -2605
rect 6833 -2639 6857 -2605
rect 6785 -2659 6857 -2639
rect 6439 -2673 6857 -2659
rect 6439 -2707 6463 -2673
rect 6497 -2707 6531 -2673
rect 6565 -2707 6731 -2673
rect 6765 -2707 6799 -2673
rect 6833 -2707 6857 -2673
rect 6439 -2731 6857 -2707
rect -941 -3157 -523 -3133
rect -941 -3191 -917 -3157
rect -883 -3191 -849 -3157
rect -815 -3191 -649 -3157
rect -615 -3191 -581 -3157
rect -547 -3191 -523 -3157
rect -941 -3205 -523 -3191
rect -941 -3225 -869 -3205
rect -941 -3259 -917 -3225
rect -883 -3259 -869 -3225
rect -941 -3425 -869 -3259
rect -595 -3225 -523 -3205
rect -595 -3259 -581 -3225
rect -547 -3259 -523 -3225
rect -941 -3459 -917 -3425
rect -883 -3459 -869 -3425
rect -941 -3479 -869 -3459
rect -595 -3425 -523 -3259
rect -595 -3459 -581 -3425
rect -547 -3459 -523 -3425
rect -595 -3479 -523 -3459
rect -941 -3493 -523 -3479
rect -941 -3527 -917 -3493
rect -883 -3527 -849 -3493
rect -815 -3527 -649 -3493
rect -615 -3527 -581 -3493
rect -547 -3527 -523 -3493
rect -941 -3551 -523 -3527
rect -121 -3157 297 -3133
rect -121 -3191 -97 -3157
rect -63 -3191 -29 -3157
rect 5 -3191 171 -3157
rect 205 -3191 239 -3157
rect 273 -3191 297 -3157
rect -121 -3205 297 -3191
rect -121 -3225 -49 -3205
rect -121 -3259 -97 -3225
rect -63 -3259 -49 -3225
rect -121 -3425 -49 -3259
rect 225 -3225 297 -3205
rect 225 -3259 239 -3225
rect 273 -3259 297 -3225
rect -121 -3459 -97 -3425
rect -63 -3459 -49 -3425
rect -121 -3479 -49 -3459
rect 225 -3425 297 -3259
rect 225 -3459 239 -3425
rect 273 -3459 297 -3425
rect 225 -3479 297 -3459
rect -121 -3493 297 -3479
rect -121 -3527 -97 -3493
rect -63 -3527 -29 -3493
rect 5 -3527 171 -3493
rect 205 -3527 239 -3493
rect 273 -3527 297 -3493
rect -121 -3551 297 -3527
rect 699 -3157 1117 -3133
rect 699 -3191 723 -3157
rect 757 -3191 791 -3157
rect 825 -3191 991 -3157
rect 1025 -3191 1059 -3157
rect 1093 -3191 1117 -3157
rect 699 -3205 1117 -3191
rect 699 -3225 771 -3205
rect 699 -3259 723 -3225
rect 757 -3259 771 -3225
rect 699 -3425 771 -3259
rect 1045 -3225 1117 -3205
rect 1045 -3259 1059 -3225
rect 1093 -3259 1117 -3225
rect 699 -3459 723 -3425
rect 757 -3459 771 -3425
rect 699 -3479 771 -3459
rect 1045 -3425 1117 -3259
rect 1045 -3459 1059 -3425
rect 1093 -3459 1117 -3425
rect 1045 -3479 1117 -3459
rect 699 -3493 1117 -3479
rect 699 -3527 723 -3493
rect 757 -3527 791 -3493
rect 825 -3527 991 -3493
rect 1025 -3527 1059 -3493
rect 1093 -3527 1117 -3493
rect 699 -3551 1117 -3527
rect 1519 -3157 1937 -3133
rect 1519 -3191 1543 -3157
rect 1577 -3191 1611 -3157
rect 1645 -3191 1811 -3157
rect 1845 -3191 1879 -3157
rect 1913 -3191 1937 -3157
rect 1519 -3205 1937 -3191
rect 1519 -3225 1591 -3205
rect 1519 -3259 1543 -3225
rect 1577 -3259 1591 -3225
rect 1519 -3425 1591 -3259
rect 1865 -3225 1937 -3205
rect 1865 -3259 1879 -3225
rect 1913 -3259 1937 -3225
rect 1519 -3459 1543 -3425
rect 1577 -3459 1591 -3425
rect 1519 -3479 1591 -3459
rect 1865 -3425 1937 -3259
rect 1865 -3459 1879 -3425
rect 1913 -3459 1937 -3425
rect 1865 -3479 1937 -3459
rect 1519 -3493 1937 -3479
rect 1519 -3527 1543 -3493
rect 1577 -3527 1611 -3493
rect 1645 -3527 1811 -3493
rect 1845 -3527 1879 -3493
rect 1913 -3527 1937 -3493
rect 1519 -3551 1937 -3527
rect 2339 -3157 2757 -3133
rect 2339 -3191 2363 -3157
rect 2397 -3191 2431 -3157
rect 2465 -3191 2631 -3157
rect 2665 -3191 2699 -3157
rect 2733 -3191 2757 -3157
rect 2339 -3205 2757 -3191
rect 2339 -3225 2411 -3205
rect 2339 -3259 2363 -3225
rect 2397 -3259 2411 -3225
rect 2339 -3425 2411 -3259
rect 2685 -3225 2757 -3205
rect 2685 -3259 2699 -3225
rect 2733 -3259 2757 -3225
rect 2339 -3459 2363 -3425
rect 2397 -3459 2411 -3425
rect 2339 -3479 2411 -3459
rect 2685 -3425 2757 -3259
rect 2685 -3459 2699 -3425
rect 2733 -3459 2757 -3425
rect 2685 -3479 2757 -3459
rect 2339 -3493 2757 -3479
rect 2339 -3527 2363 -3493
rect 2397 -3527 2431 -3493
rect 2465 -3527 2631 -3493
rect 2665 -3527 2699 -3493
rect 2733 -3527 2757 -3493
rect 2339 -3551 2757 -3527
rect 3159 -3157 3577 -3133
rect 3159 -3191 3183 -3157
rect 3217 -3191 3251 -3157
rect 3285 -3191 3451 -3157
rect 3485 -3191 3519 -3157
rect 3553 -3191 3577 -3157
rect 3159 -3205 3577 -3191
rect 3159 -3225 3231 -3205
rect 3159 -3259 3183 -3225
rect 3217 -3259 3231 -3225
rect 3159 -3425 3231 -3259
rect 3505 -3225 3577 -3205
rect 3505 -3259 3519 -3225
rect 3553 -3259 3577 -3225
rect 3159 -3459 3183 -3425
rect 3217 -3459 3231 -3425
rect 3159 -3479 3231 -3459
rect 3505 -3425 3577 -3259
rect 3505 -3459 3519 -3425
rect 3553 -3459 3577 -3425
rect 3505 -3479 3577 -3459
rect 3159 -3493 3577 -3479
rect 3159 -3527 3183 -3493
rect 3217 -3527 3251 -3493
rect 3285 -3527 3451 -3493
rect 3485 -3527 3519 -3493
rect 3553 -3527 3577 -3493
rect 3159 -3551 3577 -3527
rect 3979 -3157 4397 -3133
rect 3979 -3191 4003 -3157
rect 4037 -3191 4071 -3157
rect 4105 -3191 4271 -3157
rect 4305 -3191 4339 -3157
rect 4373 -3191 4397 -3157
rect 3979 -3205 4397 -3191
rect 3979 -3225 4051 -3205
rect 3979 -3259 4003 -3225
rect 4037 -3259 4051 -3225
rect 3979 -3425 4051 -3259
rect 4325 -3225 4397 -3205
rect 4325 -3259 4339 -3225
rect 4373 -3259 4397 -3225
rect 3979 -3459 4003 -3425
rect 4037 -3459 4051 -3425
rect 3979 -3479 4051 -3459
rect 4325 -3425 4397 -3259
rect 4325 -3459 4339 -3425
rect 4373 -3459 4397 -3425
rect 4325 -3479 4397 -3459
rect 3979 -3493 4397 -3479
rect 3979 -3527 4003 -3493
rect 4037 -3527 4071 -3493
rect 4105 -3527 4271 -3493
rect 4305 -3527 4339 -3493
rect 4373 -3527 4397 -3493
rect 3979 -3551 4397 -3527
rect 4799 -3157 5217 -3133
rect 4799 -3191 4823 -3157
rect 4857 -3191 4891 -3157
rect 4925 -3191 5091 -3157
rect 5125 -3191 5159 -3157
rect 5193 -3191 5217 -3157
rect 4799 -3205 5217 -3191
rect 4799 -3225 4871 -3205
rect 4799 -3259 4823 -3225
rect 4857 -3259 4871 -3225
rect 4799 -3425 4871 -3259
rect 5145 -3225 5217 -3205
rect 5145 -3259 5159 -3225
rect 5193 -3259 5217 -3225
rect 4799 -3459 4823 -3425
rect 4857 -3459 4871 -3425
rect 4799 -3479 4871 -3459
rect 5145 -3425 5217 -3259
rect 5145 -3459 5159 -3425
rect 5193 -3459 5217 -3425
rect 5145 -3479 5217 -3459
rect 4799 -3493 5217 -3479
rect 4799 -3527 4823 -3493
rect 4857 -3527 4891 -3493
rect 4925 -3527 5091 -3493
rect 5125 -3527 5159 -3493
rect 5193 -3527 5217 -3493
rect 4799 -3551 5217 -3527
rect 5619 -3157 6037 -3133
rect 5619 -3191 5643 -3157
rect 5677 -3191 5711 -3157
rect 5745 -3191 5911 -3157
rect 5945 -3191 5979 -3157
rect 6013 -3191 6037 -3157
rect 5619 -3205 6037 -3191
rect 5619 -3225 5691 -3205
rect 5619 -3259 5643 -3225
rect 5677 -3259 5691 -3225
rect 5619 -3425 5691 -3259
rect 5965 -3225 6037 -3205
rect 5965 -3259 5979 -3225
rect 6013 -3259 6037 -3225
rect 5619 -3459 5643 -3425
rect 5677 -3459 5691 -3425
rect 5619 -3479 5691 -3459
rect 5965 -3425 6037 -3259
rect 5965 -3459 5979 -3425
rect 6013 -3459 6037 -3425
rect 5965 -3479 6037 -3459
rect 5619 -3493 6037 -3479
rect 5619 -3527 5643 -3493
rect 5677 -3527 5711 -3493
rect 5745 -3527 5911 -3493
rect 5945 -3527 5979 -3493
rect 6013 -3527 6037 -3493
rect 5619 -3551 6037 -3527
rect 6439 -3157 6857 -3133
rect 6439 -3191 6463 -3157
rect 6497 -3191 6531 -3157
rect 6565 -3191 6731 -3157
rect 6765 -3191 6799 -3157
rect 6833 -3191 6857 -3157
rect 6439 -3205 6857 -3191
rect 6439 -3225 6511 -3205
rect 6439 -3259 6463 -3225
rect 6497 -3259 6511 -3225
rect 6439 -3425 6511 -3259
rect 6785 -3225 6857 -3205
rect 6785 -3259 6799 -3225
rect 6833 -3259 6857 -3225
rect 6439 -3459 6463 -3425
rect 6497 -3459 6511 -3425
rect 6439 -3479 6511 -3459
rect 6785 -3425 6857 -3259
rect 6785 -3459 6799 -3425
rect 6833 -3459 6857 -3425
rect 6785 -3479 6857 -3459
rect 6439 -3493 6857 -3479
rect 6439 -3527 6463 -3493
rect 6497 -3527 6531 -3493
rect 6565 -3527 6731 -3493
rect 6765 -3527 6799 -3493
rect 6833 -3527 6857 -3493
rect 6439 -3551 6857 -3527
rect -941 -3977 -523 -3953
rect -941 -4011 -917 -3977
rect -883 -4011 -849 -3977
rect -815 -4011 -649 -3977
rect -615 -4011 -581 -3977
rect -547 -4011 -523 -3977
rect -941 -4025 -523 -4011
rect -941 -4045 -869 -4025
rect -941 -4079 -917 -4045
rect -883 -4079 -869 -4045
rect -941 -4245 -869 -4079
rect -595 -4045 -523 -4025
rect -595 -4079 -581 -4045
rect -547 -4079 -523 -4045
rect -941 -4279 -917 -4245
rect -883 -4279 -869 -4245
rect -941 -4299 -869 -4279
rect -595 -4245 -523 -4079
rect -595 -4279 -581 -4245
rect -547 -4279 -523 -4245
rect -595 -4299 -523 -4279
rect -941 -4313 -523 -4299
rect -941 -4347 -917 -4313
rect -883 -4347 -849 -4313
rect -815 -4347 -649 -4313
rect -615 -4347 -581 -4313
rect -547 -4347 -523 -4313
rect -941 -4371 -523 -4347
rect -121 -3977 297 -3953
rect -121 -4011 -97 -3977
rect -63 -4011 -29 -3977
rect 5 -4011 171 -3977
rect 205 -4011 239 -3977
rect 273 -4011 297 -3977
rect -121 -4025 297 -4011
rect -121 -4045 -49 -4025
rect -121 -4079 -97 -4045
rect -63 -4079 -49 -4045
rect -121 -4245 -49 -4079
rect 225 -4045 297 -4025
rect 225 -4079 239 -4045
rect 273 -4079 297 -4045
rect -121 -4279 -97 -4245
rect -63 -4279 -49 -4245
rect -121 -4299 -49 -4279
rect 225 -4245 297 -4079
rect 225 -4279 239 -4245
rect 273 -4279 297 -4245
rect 225 -4299 297 -4279
rect -121 -4313 297 -4299
rect -121 -4347 -97 -4313
rect -63 -4347 -29 -4313
rect 5 -4347 171 -4313
rect 205 -4347 239 -4313
rect 273 -4347 297 -4313
rect -121 -4371 297 -4347
rect 699 -3977 1117 -3953
rect 699 -4011 723 -3977
rect 757 -4011 791 -3977
rect 825 -4011 991 -3977
rect 1025 -4011 1059 -3977
rect 1093 -4011 1117 -3977
rect 699 -4025 1117 -4011
rect 699 -4045 771 -4025
rect 699 -4079 723 -4045
rect 757 -4079 771 -4045
rect 699 -4245 771 -4079
rect 1045 -4045 1117 -4025
rect 1045 -4079 1059 -4045
rect 1093 -4079 1117 -4045
rect 699 -4279 723 -4245
rect 757 -4279 771 -4245
rect 699 -4299 771 -4279
rect 1045 -4245 1117 -4079
rect 1045 -4279 1059 -4245
rect 1093 -4279 1117 -4245
rect 1045 -4299 1117 -4279
rect 699 -4313 1117 -4299
rect 699 -4347 723 -4313
rect 757 -4347 791 -4313
rect 825 -4347 991 -4313
rect 1025 -4347 1059 -4313
rect 1093 -4347 1117 -4313
rect 699 -4371 1117 -4347
rect 1519 -3977 1937 -3953
rect 1519 -4011 1543 -3977
rect 1577 -4011 1611 -3977
rect 1645 -4011 1811 -3977
rect 1845 -4011 1879 -3977
rect 1913 -4011 1937 -3977
rect 1519 -4025 1937 -4011
rect 1519 -4045 1591 -4025
rect 1519 -4079 1543 -4045
rect 1577 -4079 1591 -4045
rect 1519 -4245 1591 -4079
rect 1865 -4045 1937 -4025
rect 1865 -4079 1879 -4045
rect 1913 -4079 1937 -4045
rect 1519 -4279 1543 -4245
rect 1577 -4279 1591 -4245
rect 1519 -4299 1591 -4279
rect 1865 -4245 1937 -4079
rect 1865 -4279 1879 -4245
rect 1913 -4279 1937 -4245
rect 1865 -4299 1937 -4279
rect 1519 -4313 1937 -4299
rect 1519 -4347 1543 -4313
rect 1577 -4347 1611 -4313
rect 1645 -4347 1811 -4313
rect 1845 -4347 1879 -4313
rect 1913 -4347 1937 -4313
rect 1519 -4371 1937 -4347
rect 2339 -3977 2757 -3953
rect 2339 -4011 2363 -3977
rect 2397 -4011 2431 -3977
rect 2465 -4011 2631 -3977
rect 2665 -4011 2699 -3977
rect 2733 -4011 2757 -3977
rect 2339 -4025 2757 -4011
rect 2339 -4045 2411 -4025
rect 2339 -4079 2363 -4045
rect 2397 -4079 2411 -4045
rect 2339 -4245 2411 -4079
rect 2685 -4045 2757 -4025
rect 2685 -4079 2699 -4045
rect 2733 -4079 2757 -4045
rect 2339 -4279 2363 -4245
rect 2397 -4279 2411 -4245
rect 2339 -4299 2411 -4279
rect 2685 -4245 2757 -4079
rect 2685 -4279 2699 -4245
rect 2733 -4279 2757 -4245
rect 2685 -4299 2757 -4279
rect 2339 -4313 2757 -4299
rect 2339 -4347 2363 -4313
rect 2397 -4347 2431 -4313
rect 2465 -4347 2631 -4313
rect 2665 -4347 2699 -4313
rect 2733 -4347 2757 -4313
rect 2339 -4371 2757 -4347
rect 3159 -3977 3577 -3953
rect 3159 -4011 3183 -3977
rect 3217 -4011 3251 -3977
rect 3285 -4011 3451 -3977
rect 3485 -4011 3519 -3977
rect 3553 -4011 3577 -3977
rect 3159 -4025 3577 -4011
rect 3159 -4045 3231 -4025
rect 3159 -4079 3183 -4045
rect 3217 -4079 3231 -4045
rect 3159 -4245 3231 -4079
rect 3505 -4045 3577 -4025
rect 3505 -4079 3519 -4045
rect 3553 -4079 3577 -4045
rect 3159 -4279 3183 -4245
rect 3217 -4279 3231 -4245
rect 3159 -4299 3231 -4279
rect 3505 -4245 3577 -4079
rect 3505 -4279 3519 -4245
rect 3553 -4279 3577 -4245
rect 3505 -4299 3577 -4279
rect 3159 -4313 3577 -4299
rect 3159 -4347 3183 -4313
rect 3217 -4347 3251 -4313
rect 3285 -4347 3451 -4313
rect 3485 -4347 3519 -4313
rect 3553 -4347 3577 -4313
rect 3159 -4371 3577 -4347
rect 3979 -3977 4397 -3953
rect 3979 -4011 4003 -3977
rect 4037 -4011 4071 -3977
rect 4105 -4011 4271 -3977
rect 4305 -4011 4339 -3977
rect 4373 -4011 4397 -3977
rect 3979 -4025 4397 -4011
rect 3979 -4045 4051 -4025
rect 3979 -4079 4003 -4045
rect 4037 -4079 4051 -4045
rect 3979 -4245 4051 -4079
rect 4325 -4045 4397 -4025
rect 4325 -4079 4339 -4045
rect 4373 -4079 4397 -4045
rect 3979 -4279 4003 -4245
rect 4037 -4279 4051 -4245
rect 3979 -4299 4051 -4279
rect 4325 -4245 4397 -4079
rect 4325 -4279 4339 -4245
rect 4373 -4279 4397 -4245
rect 4325 -4299 4397 -4279
rect 3979 -4313 4397 -4299
rect 3979 -4347 4003 -4313
rect 4037 -4347 4071 -4313
rect 4105 -4347 4271 -4313
rect 4305 -4347 4339 -4313
rect 4373 -4347 4397 -4313
rect 3979 -4371 4397 -4347
rect 4799 -3977 5217 -3953
rect 4799 -4011 4823 -3977
rect 4857 -4011 4891 -3977
rect 4925 -4011 5091 -3977
rect 5125 -4011 5159 -3977
rect 5193 -4011 5217 -3977
rect 4799 -4025 5217 -4011
rect 4799 -4045 4871 -4025
rect 4799 -4079 4823 -4045
rect 4857 -4079 4871 -4045
rect 4799 -4245 4871 -4079
rect 5145 -4045 5217 -4025
rect 5145 -4079 5159 -4045
rect 5193 -4079 5217 -4045
rect 4799 -4279 4823 -4245
rect 4857 -4279 4871 -4245
rect 4799 -4299 4871 -4279
rect 5145 -4245 5217 -4079
rect 5145 -4279 5159 -4245
rect 5193 -4279 5217 -4245
rect 5145 -4299 5217 -4279
rect 4799 -4313 5217 -4299
rect 4799 -4347 4823 -4313
rect 4857 -4347 4891 -4313
rect 4925 -4347 5091 -4313
rect 5125 -4347 5159 -4313
rect 5193 -4347 5217 -4313
rect 4799 -4371 5217 -4347
rect 5619 -3977 6037 -3953
rect 5619 -4011 5643 -3977
rect 5677 -4011 5711 -3977
rect 5745 -4011 5911 -3977
rect 5945 -4011 5979 -3977
rect 6013 -4011 6037 -3977
rect 5619 -4025 6037 -4011
rect 5619 -4045 5691 -4025
rect 5619 -4079 5643 -4045
rect 5677 -4079 5691 -4045
rect 5619 -4245 5691 -4079
rect 5965 -4045 6037 -4025
rect 5965 -4079 5979 -4045
rect 6013 -4079 6037 -4045
rect 5619 -4279 5643 -4245
rect 5677 -4279 5691 -4245
rect 5619 -4299 5691 -4279
rect 5965 -4245 6037 -4079
rect 5965 -4279 5979 -4245
rect 6013 -4279 6037 -4245
rect 5965 -4299 6037 -4279
rect 5619 -4313 6037 -4299
rect 5619 -4347 5643 -4313
rect 5677 -4347 5711 -4313
rect 5745 -4347 5911 -4313
rect 5945 -4347 5979 -4313
rect 6013 -4347 6037 -4313
rect 5619 -4371 6037 -4347
rect 6439 -3977 6857 -3953
rect 6439 -4011 6463 -3977
rect 6497 -4011 6531 -3977
rect 6565 -4011 6731 -3977
rect 6765 -4011 6799 -3977
rect 6833 -4011 6857 -3977
rect 6439 -4025 6857 -4011
rect 6439 -4045 6511 -4025
rect 6439 -4079 6463 -4045
rect 6497 -4079 6511 -4045
rect 6439 -4245 6511 -4079
rect 6785 -4045 6857 -4025
rect 6785 -4079 6799 -4045
rect 6833 -4079 6857 -4045
rect 6439 -4279 6463 -4245
rect 6497 -4279 6511 -4245
rect 6439 -4299 6511 -4279
rect 6785 -4245 6857 -4079
rect 6785 -4279 6799 -4245
rect 6833 -4279 6857 -4245
rect 6785 -4299 6857 -4279
rect 6439 -4313 6857 -4299
rect 6439 -4347 6463 -4313
rect 6497 -4347 6531 -4313
rect 6565 -4347 6731 -4313
rect 6765 -4347 6799 -4313
rect 6833 -4347 6857 -4313
rect 6439 -4371 6857 -4347
<< psubdiffcont >>
rect -1070 -578 -1036 -544
rect -1002 -578 -968 -544
rect -934 -578 -900 -544
rect -866 -578 -832 -544
rect -632 -578 -598 -544
rect -564 -578 -530 -544
rect -496 -578 -462 -544
rect -428 -578 -394 -544
rect -1070 -646 -1036 -612
rect -428 -646 -394 -612
rect -1070 -714 -1036 -680
rect -1070 -782 -1036 -748
rect -1070 -1016 -1036 -982
rect -1070 -1084 -1036 -1050
rect -428 -714 -394 -680
rect -428 -782 -394 -748
rect -428 -1016 -394 -982
rect -428 -1084 -394 -1050
rect -1070 -1152 -1036 -1118
rect -428 -1152 -394 -1118
rect -1070 -1220 -1036 -1186
rect -1002 -1220 -968 -1186
rect -934 -1220 -900 -1186
rect -866 -1220 -832 -1186
rect -632 -1220 -598 -1186
rect -564 -1220 -530 -1186
rect -496 -1220 -462 -1186
rect -428 -1220 -394 -1186
rect -250 -578 -216 -544
rect -182 -578 -148 -544
rect -114 -578 -80 -544
rect -46 -578 -12 -544
rect 188 -578 222 -544
rect 256 -578 290 -544
rect 324 -578 358 -544
rect 392 -578 426 -544
rect -250 -646 -216 -612
rect 392 -646 426 -612
rect -250 -714 -216 -680
rect -250 -782 -216 -748
rect -250 -1016 -216 -982
rect -250 -1084 -216 -1050
rect 392 -714 426 -680
rect 392 -782 426 -748
rect 392 -1016 426 -982
rect 392 -1084 426 -1050
rect -250 -1152 -216 -1118
rect 392 -1152 426 -1118
rect -250 -1220 -216 -1186
rect -182 -1220 -148 -1186
rect -114 -1220 -80 -1186
rect -46 -1220 -12 -1186
rect 188 -1220 222 -1186
rect 256 -1220 290 -1186
rect 324 -1220 358 -1186
rect 392 -1220 426 -1186
rect 570 -578 604 -544
rect 638 -578 672 -544
rect 706 -578 740 -544
rect 774 -578 808 -544
rect 1008 -578 1042 -544
rect 1076 -578 1110 -544
rect 1144 -578 1178 -544
rect 1212 -578 1246 -544
rect 570 -646 604 -612
rect 1212 -646 1246 -612
rect 570 -714 604 -680
rect 570 -782 604 -748
rect 570 -1016 604 -982
rect 570 -1084 604 -1050
rect 1212 -714 1246 -680
rect 1212 -782 1246 -748
rect 1212 -1016 1246 -982
rect 1212 -1084 1246 -1050
rect 570 -1152 604 -1118
rect 1212 -1152 1246 -1118
rect 570 -1220 604 -1186
rect 638 -1220 672 -1186
rect 706 -1220 740 -1186
rect 774 -1220 808 -1186
rect 1008 -1220 1042 -1186
rect 1076 -1220 1110 -1186
rect 1144 -1220 1178 -1186
rect 1212 -1220 1246 -1186
rect 1390 -578 1424 -544
rect 1458 -578 1492 -544
rect 1526 -578 1560 -544
rect 1594 -578 1628 -544
rect 1828 -578 1862 -544
rect 1896 -578 1930 -544
rect 1964 -578 1998 -544
rect 2032 -578 2066 -544
rect 1390 -646 1424 -612
rect 2032 -646 2066 -612
rect 1390 -714 1424 -680
rect 1390 -782 1424 -748
rect 1390 -1016 1424 -982
rect 1390 -1084 1424 -1050
rect 2032 -714 2066 -680
rect 2032 -782 2066 -748
rect 2032 -1016 2066 -982
rect 2032 -1084 2066 -1050
rect 1390 -1152 1424 -1118
rect 2032 -1152 2066 -1118
rect 1390 -1220 1424 -1186
rect 1458 -1220 1492 -1186
rect 1526 -1220 1560 -1186
rect 1594 -1220 1628 -1186
rect 1828 -1220 1862 -1186
rect 1896 -1220 1930 -1186
rect 1964 -1220 1998 -1186
rect 2032 -1220 2066 -1186
rect 2210 -578 2244 -544
rect 2278 -578 2312 -544
rect 2346 -578 2380 -544
rect 2414 -578 2448 -544
rect 2648 -578 2682 -544
rect 2716 -578 2750 -544
rect 2784 -578 2818 -544
rect 2852 -578 2886 -544
rect 2210 -646 2244 -612
rect 2852 -646 2886 -612
rect 2210 -714 2244 -680
rect 2210 -782 2244 -748
rect 2210 -1016 2244 -982
rect 2210 -1084 2244 -1050
rect 2852 -714 2886 -680
rect 2852 -782 2886 -748
rect 2852 -1016 2886 -982
rect 2852 -1084 2886 -1050
rect 2210 -1152 2244 -1118
rect 2852 -1152 2886 -1118
rect 2210 -1220 2244 -1186
rect 2278 -1220 2312 -1186
rect 2346 -1220 2380 -1186
rect 2414 -1220 2448 -1186
rect 2648 -1220 2682 -1186
rect 2716 -1220 2750 -1186
rect 2784 -1220 2818 -1186
rect 2852 -1220 2886 -1186
rect 3030 -578 3064 -544
rect 3098 -578 3132 -544
rect 3166 -578 3200 -544
rect 3234 -578 3268 -544
rect 3468 -578 3502 -544
rect 3536 -578 3570 -544
rect 3604 -578 3638 -544
rect 3672 -578 3706 -544
rect 3030 -646 3064 -612
rect 3672 -646 3706 -612
rect 3030 -714 3064 -680
rect 3030 -782 3064 -748
rect 3030 -1016 3064 -982
rect 3030 -1084 3064 -1050
rect 3672 -714 3706 -680
rect 3672 -782 3706 -748
rect 3672 -1016 3706 -982
rect 3672 -1084 3706 -1050
rect 3030 -1152 3064 -1118
rect 3672 -1152 3706 -1118
rect 3030 -1220 3064 -1186
rect 3098 -1220 3132 -1186
rect 3166 -1220 3200 -1186
rect 3234 -1220 3268 -1186
rect 3468 -1220 3502 -1186
rect 3536 -1220 3570 -1186
rect 3604 -1220 3638 -1186
rect 3672 -1220 3706 -1186
rect 3850 -578 3884 -544
rect 3918 -578 3952 -544
rect 3986 -578 4020 -544
rect 4054 -578 4088 -544
rect 4288 -578 4322 -544
rect 4356 -578 4390 -544
rect 4424 -578 4458 -544
rect 4492 -578 4526 -544
rect 3850 -646 3884 -612
rect 4492 -646 4526 -612
rect 3850 -714 3884 -680
rect 3850 -782 3884 -748
rect 3850 -1016 3884 -982
rect 3850 -1084 3884 -1050
rect 4492 -714 4526 -680
rect 4492 -782 4526 -748
rect 4492 -1016 4526 -982
rect 4492 -1084 4526 -1050
rect 3850 -1152 3884 -1118
rect 4492 -1152 4526 -1118
rect 3850 -1220 3884 -1186
rect 3918 -1220 3952 -1186
rect 3986 -1220 4020 -1186
rect 4054 -1220 4088 -1186
rect 4288 -1220 4322 -1186
rect 4356 -1220 4390 -1186
rect 4424 -1220 4458 -1186
rect 4492 -1220 4526 -1186
rect 4670 -578 4704 -544
rect 4738 -578 4772 -544
rect 4806 -578 4840 -544
rect 4874 -578 4908 -544
rect 5108 -578 5142 -544
rect 5176 -578 5210 -544
rect 5244 -578 5278 -544
rect 5312 -578 5346 -544
rect 4670 -646 4704 -612
rect 5312 -646 5346 -612
rect 4670 -714 4704 -680
rect 4670 -782 4704 -748
rect 4670 -1016 4704 -982
rect 4670 -1084 4704 -1050
rect 5312 -714 5346 -680
rect 5312 -782 5346 -748
rect 5312 -1016 5346 -982
rect 5312 -1084 5346 -1050
rect 4670 -1152 4704 -1118
rect 5312 -1152 5346 -1118
rect 4670 -1220 4704 -1186
rect 4738 -1220 4772 -1186
rect 4806 -1220 4840 -1186
rect 4874 -1220 4908 -1186
rect 5108 -1220 5142 -1186
rect 5176 -1220 5210 -1186
rect 5244 -1220 5278 -1186
rect 5312 -1220 5346 -1186
rect 5490 -578 5524 -544
rect 5558 -578 5592 -544
rect 5626 -578 5660 -544
rect 5694 -578 5728 -544
rect 5928 -578 5962 -544
rect 5996 -578 6030 -544
rect 6064 -578 6098 -544
rect 6132 -578 6166 -544
rect 5490 -646 5524 -612
rect 6132 -646 6166 -612
rect 5490 -714 5524 -680
rect 5490 -782 5524 -748
rect 5490 -1016 5524 -982
rect 5490 -1084 5524 -1050
rect 6132 -714 6166 -680
rect 6132 -782 6166 -748
rect 6132 -1016 6166 -982
rect 6132 -1084 6166 -1050
rect 5490 -1152 5524 -1118
rect 6132 -1152 6166 -1118
rect 5490 -1220 5524 -1186
rect 5558 -1220 5592 -1186
rect 5626 -1220 5660 -1186
rect 5694 -1220 5728 -1186
rect 5928 -1220 5962 -1186
rect 5996 -1220 6030 -1186
rect 6064 -1220 6098 -1186
rect 6132 -1220 6166 -1186
rect 6310 -578 6344 -544
rect 6378 -578 6412 -544
rect 6446 -578 6480 -544
rect 6514 -578 6548 -544
rect 6748 -578 6782 -544
rect 6816 -578 6850 -544
rect 6884 -578 6918 -544
rect 6952 -578 6986 -544
rect 6310 -646 6344 -612
rect 6952 -646 6986 -612
rect 6310 -714 6344 -680
rect 6310 -782 6344 -748
rect 6310 -1016 6344 -982
rect 6310 -1084 6344 -1050
rect 6952 -714 6986 -680
rect 6952 -782 6986 -748
rect 6952 -1016 6986 -982
rect 6952 -1084 6986 -1050
rect 6310 -1152 6344 -1118
rect 6952 -1152 6986 -1118
rect 6310 -1220 6344 -1186
rect 6378 -1220 6412 -1186
rect 6446 -1220 6480 -1186
rect 6514 -1220 6548 -1186
rect 6748 -1220 6782 -1186
rect 6816 -1220 6850 -1186
rect 6884 -1220 6918 -1186
rect 6952 -1220 6986 -1186
rect 7160 -578 7194 -544
rect 7228 -578 7262 -544
rect 7296 -578 7330 -544
rect 7364 -578 7398 -544
rect 7598 -578 7632 -544
rect 7666 -578 7700 -544
rect 7734 -578 7768 -544
rect 7802 -578 7836 -544
rect 7160 -646 7194 -612
rect 7802 -646 7836 -612
rect 7160 -714 7194 -680
rect 7160 -782 7194 -748
rect 7160 -1016 7194 -982
rect 7160 -1084 7194 -1050
rect 7802 -714 7836 -680
rect 7802 -782 7836 -748
rect 7802 -1016 7836 -982
rect 7802 -1084 7836 -1050
rect 7160 -1152 7194 -1118
rect 7802 -1152 7836 -1118
rect 7160 -1220 7194 -1186
rect 7228 -1220 7262 -1186
rect 7296 -1220 7330 -1186
rect 7364 -1220 7398 -1186
rect 7598 -1220 7632 -1186
rect 7666 -1220 7700 -1186
rect 7734 -1220 7768 -1186
rect 7802 -1220 7836 -1186
rect -1070 -1398 -1036 -1364
rect -1002 -1398 -968 -1364
rect -934 -1398 -900 -1364
rect -866 -1398 -832 -1364
rect -632 -1398 -598 -1364
rect -564 -1398 -530 -1364
rect -496 -1398 -462 -1364
rect -428 -1398 -394 -1364
rect -1070 -1466 -1036 -1432
rect -428 -1466 -394 -1432
rect -1070 -1534 -1036 -1500
rect -1070 -1602 -1036 -1568
rect -1070 -1836 -1036 -1802
rect -1070 -1904 -1036 -1870
rect -428 -1534 -394 -1500
rect -428 -1602 -394 -1568
rect -428 -1836 -394 -1802
rect -428 -1904 -394 -1870
rect -1070 -1972 -1036 -1938
rect -428 -1972 -394 -1938
rect -1070 -2040 -1036 -2006
rect -1002 -2040 -968 -2006
rect -934 -2040 -900 -2006
rect -866 -2040 -832 -2006
rect -632 -2040 -598 -2006
rect -564 -2040 -530 -2006
rect -496 -2040 -462 -2006
rect -428 -2040 -394 -2006
rect -250 -1398 -216 -1364
rect -182 -1398 -148 -1364
rect -114 -1398 -80 -1364
rect -46 -1398 -12 -1364
rect 188 -1398 222 -1364
rect 256 -1398 290 -1364
rect 324 -1398 358 -1364
rect 392 -1398 426 -1364
rect -250 -1466 -216 -1432
rect 392 -1466 426 -1432
rect -250 -1534 -216 -1500
rect -250 -1602 -216 -1568
rect -250 -1836 -216 -1802
rect -250 -1904 -216 -1870
rect 392 -1534 426 -1500
rect 392 -1602 426 -1568
rect 392 -1836 426 -1802
rect 392 -1904 426 -1870
rect -250 -1972 -216 -1938
rect 392 -1972 426 -1938
rect -250 -2040 -216 -2006
rect -182 -2040 -148 -2006
rect -114 -2040 -80 -2006
rect -46 -2040 -12 -2006
rect 188 -2040 222 -2006
rect 256 -2040 290 -2006
rect 324 -2040 358 -2006
rect 392 -2040 426 -2006
rect 570 -1398 604 -1364
rect 638 -1398 672 -1364
rect 706 -1398 740 -1364
rect 774 -1398 808 -1364
rect 1008 -1398 1042 -1364
rect 1076 -1398 1110 -1364
rect 1144 -1398 1178 -1364
rect 1212 -1398 1246 -1364
rect 570 -1466 604 -1432
rect 1212 -1466 1246 -1432
rect 570 -1534 604 -1500
rect 570 -1602 604 -1568
rect 570 -1836 604 -1802
rect 570 -1904 604 -1870
rect 1212 -1534 1246 -1500
rect 1212 -1602 1246 -1568
rect 1212 -1836 1246 -1802
rect 1212 -1904 1246 -1870
rect 570 -1972 604 -1938
rect 1212 -1972 1246 -1938
rect 570 -2040 604 -2006
rect 638 -2040 672 -2006
rect 706 -2040 740 -2006
rect 774 -2040 808 -2006
rect 1008 -2040 1042 -2006
rect 1076 -2040 1110 -2006
rect 1144 -2040 1178 -2006
rect 1212 -2040 1246 -2006
rect 1390 -1398 1424 -1364
rect 1458 -1398 1492 -1364
rect 1526 -1398 1560 -1364
rect 1594 -1398 1628 -1364
rect 1828 -1398 1862 -1364
rect 1896 -1398 1930 -1364
rect 1964 -1398 1998 -1364
rect 2032 -1398 2066 -1364
rect 1390 -1466 1424 -1432
rect 2032 -1466 2066 -1432
rect 1390 -1534 1424 -1500
rect 1390 -1602 1424 -1568
rect 1390 -1836 1424 -1802
rect 1390 -1904 1424 -1870
rect 2032 -1534 2066 -1500
rect 2032 -1602 2066 -1568
rect 2032 -1836 2066 -1802
rect 2032 -1904 2066 -1870
rect 1390 -1972 1424 -1938
rect 2032 -1972 2066 -1938
rect 1390 -2040 1424 -2006
rect 1458 -2040 1492 -2006
rect 1526 -2040 1560 -2006
rect 1594 -2040 1628 -2006
rect 1828 -2040 1862 -2006
rect 1896 -2040 1930 -2006
rect 1964 -2040 1998 -2006
rect 2032 -2040 2066 -2006
rect 2210 -1398 2244 -1364
rect 2278 -1398 2312 -1364
rect 2346 -1398 2380 -1364
rect 2414 -1398 2448 -1364
rect 2648 -1398 2682 -1364
rect 2716 -1398 2750 -1364
rect 2784 -1398 2818 -1364
rect 2852 -1398 2886 -1364
rect 2210 -1466 2244 -1432
rect 2852 -1466 2886 -1432
rect 2210 -1534 2244 -1500
rect 2210 -1602 2244 -1568
rect 2210 -1836 2244 -1802
rect 2210 -1904 2244 -1870
rect 2852 -1534 2886 -1500
rect 2852 -1602 2886 -1568
rect 2852 -1836 2886 -1802
rect 2852 -1904 2886 -1870
rect 2210 -1972 2244 -1938
rect 2852 -1972 2886 -1938
rect 2210 -2040 2244 -2006
rect 2278 -2040 2312 -2006
rect 2346 -2040 2380 -2006
rect 2414 -2040 2448 -2006
rect 2648 -2040 2682 -2006
rect 2716 -2040 2750 -2006
rect 2784 -2040 2818 -2006
rect 2852 -2040 2886 -2006
rect 3030 -1398 3064 -1364
rect 3098 -1398 3132 -1364
rect 3166 -1398 3200 -1364
rect 3234 -1398 3268 -1364
rect 3468 -1398 3502 -1364
rect 3536 -1398 3570 -1364
rect 3604 -1398 3638 -1364
rect 3672 -1398 3706 -1364
rect 3030 -1466 3064 -1432
rect 3672 -1466 3706 -1432
rect 3030 -1534 3064 -1500
rect 3030 -1602 3064 -1568
rect 3030 -1836 3064 -1802
rect 3030 -1904 3064 -1870
rect 3672 -1534 3706 -1500
rect 3672 -1602 3706 -1568
rect 3672 -1836 3706 -1802
rect 3672 -1904 3706 -1870
rect 3030 -1972 3064 -1938
rect 3672 -1972 3706 -1938
rect 3030 -2040 3064 -2006
rect 3098 -2040 3132 -2006
rect 3166 -2040 3200 -2006
rect 3234 -2040 3268 -2006
rect 3468 -2040 3502 -2006
rect 3536 -2040 3570 -2006
rect 3604 -2040 3638 -2006
rect 3672 -2040 3706 -2006
rect 3850 -1398 3884 -1364
rect 3918 -1398 3952 -1364
rect 3986 -1398 4020 -1364
rect 4054 -1398 4088 -1364
rect 4288 -1398 4322 -1364
rect 4356 -1398 4390 -1364
rect 4424 -1398 4458 -1364
rect 4492 -1398 4526 -1364
rect 3850 -1466 3884 -1432
rect 4492 -1466 4526 -1432
rect 3850 -1534 3884 -1500
rect 3850 -1602 3884 -1568
rect 3850 -1836 3884 -1802
rect 3850 -1904 3884 -1870
rect 4492 -1534 4526 -1500
rect 4492 -1602 4526 -1568
rect 4492 -1836 4526 -1802
rect 4492 -1904 4526 -1870
rect 3850 -1972 3884 -1938
rect 4492 -1972 4526 -1938
rect 3850 -2040 3884 -2006
rect 3918 -2040 3952 -2006
rect 3986 -2040 4020 -2006
rect 4054 -2040 4088 -2006
rect 4288 -2040 4322 -2006
rect 4356 -2040 4390 -2006
rect 4424 -2040 4458 -2006
rect 4492 -2040 4526 -2006
rect 4670 -1398 4704 -1364
rect 4738 -1398 4772 -1364
rect 4806 -1398 4840 -1364
rect 4874 -1398 4908 -1364
rect 5108 -1398 5142 -1364
rect 5176 -1398 5210 -1364
rect 5244 -1398 5278 -1364
rect 5312 -1398 5346 -1364
rect 4670 -1466 4704 -1432
rect 5312 -1466 5346 -1432
rect 4670 -1534 4704 -1500
rect 4670 -1602 4704 -1568
rect 4670 -1836 4704 -1802
rect 4670 -1904 4704 -1870
rect 5312 -1534 5346 -1500
rect 5312 -1602 5346 -1568
rect 5312 -1836 5346 -1802
rect 5312 -1904 5346 -1870
rect 4670 -1972 4704 -1938
rect 5312 -1972 5346 -1938
rect 4670 -2040 4704 -2006
rect 4738 -2040 4772 -2006
rect 4806 -2040 4840 -2006
rect 4874 -2040 4908 -2006
rect 5108 -2040 5142 -2006
rect 5176 -2040 5210 -2006
rect 5244 -2040 5278 -2006
rect 5312 -2040 5346 -2006
rect 5490 -1398 5524 -1364
rect 5558 -1398 5592 -1364
rect 5626 -1398 5660 -1364
rect 5694 -1398 5728 -1364
rect 5928 -1398 5962 -1364
rect 5996 -1398 6030 -1364
rect 6064 -1398 6098 -1364
rect 6132 -1398 6166 -1364
rect 5490 -1466 5524 -1432
rect 6132 -1466 6166 -1432
rect 5490 -1534 5524 -1500
rect 5490 -1602 5524 -1568
rect 5490 -1836 5524 -1802
rect 5490 -1904 5524 -1870
rect 6132 -1534 6166 -1500
rect 6132 -1602 6166 -1568
rect 6132 -1836 6166 -1802
rect 6132 -1904 6166 -1870
rect 5490 -1972 5524 -1938
rect 6132 -1972 6166 -1938
rect 5490 -2040 5524 -2006
rect 5558 -2040 5592 -2006
rect 5626 -2040 5660 -2006
rect 5694 -2040 5728 -2006
rect 5928 -2040 5962 -2006
rect 5996 -2040 6030 -2006
rect 6064 -2040 6098 -2006
rect 6132 -2040 6166 -2006
rect 6310 -1398 6344 -1364
rect 6378 -1398 6412 -1364
rect 6446 -1398 6480 -1364
rect 6514 -1398 6548 -1364
rect 6748 -1398 6782 -1364
rect 6816 -1398 6850 -1364
rect 6884 -1398 6918 -1364
rect 6952 -1398 6986 -1364
rect 6310 -1466 6344 -1432
rect 6952 -1466 6986 -1432
rect 6310 -1534 6344 -1500
rect 6310 -1602 6344 -1568
rect 6310 -1836 6344 -1802
rect 6310 -1904 6344 -1870
rect 6952 -1534 6986 -1500
rect 6952 -1602 6986 -1568
rect 6952 -1836 6986 -1802
rect 6952 -1904 6986 -1870
rect 6310 -1972 6344 -1938
rect 6952 -1972 6986 -1938
rect 6310 -2040 6344 -2006
rect 6378 -2040 6412 -2006
rect 6446 -2040 6480 -2006
rect 6514 -2040 6548 -2006
rect 6748 -2040 6782 -2006
rect 6816 -2040 6850 -2006
rect 6884 -2040 6918 -2006
rect 6952 -2040 6986 -2006
rect -1070 -2218 -1036 -2184
rect -1002 -2218 -968 -2184
rect -934 -2218 -900 -2184
rect -866 -2218 -832 -2184
rect -632 -2218 -598 -2184
rect -564 -2218 -530 -2184
rect -496 -2218 -462 -2184
rect -428 -2218 -394 -2184
rect -1070 -2286 -1036 -2252
rect -428 -2286 -394 -2252
rect -1070 -2354 -1036 -2320
rect -1070 -2422 -1036 -2388
rect -1070 -2656 -1036 -2622
rect -1070 -2724 -1036 -2690
rect -428 -2354 -394 -2320
rect -428 -2422 -394 -2388
rect -428 -2656 -394 -2622
rect -428 -2724 -394 -2690
rect -1070 -2792 -1036 -2758
rect -428 -2792 -394 -2758
rect -1070 -2860 -1036 -2826
rect -1002 -2860 -968 -2826
rect -934 -2860 -900 -2826
rect -866 -2860 -832 -2826
rect -632 -2860 -598 -2826
rect -564 -2860 -530 -2826
rect -496 -2860 -462 -2826
rect -428 -2860 -394 -2826
rect -250 -2218 -216 -2184
rect -182 -2218 -148 -2184
rect -114 -2218 -80 -2184
rect -46 -2218 -12 -2184
rect 188 -2218 222 -2184
rect 256 -2218 290 -2184
rect 324 -2218 358 -2184
rect 392 -2218 426 -2184
rect -250 -2286 -216 -2252
rect 392 -2286 426 -2252
rect -250 -2354 -216 -2320
rect -250 -2422 -216 -2388
rect -250 -2656 -216 -2622
rect -250 -2724 -216 -2690
rect 392 -2354 426 -2320
rect 392 -2422 426 -2388
rect 392 -2656 426 -2622
rect 392 -2724 426 -2690
rect -250 -2792 -216 -2758
rect 392 -2792 426 -2758
rect -250 -2860 -216 -2826
rect -182 -2860 -148 -2826
rect -114 -2860 -80 -2826
rect -46 -2860 -12 -2826
rect 188 -2860 222 -2826
rect 256 -2860 290 -2826
rect 324 -2860 358 -2826
rect 392 -2860 426 -2826
rect 570 -2218 604 -2184
rect 638 -2218 672 -2184
rect 706 -2218 740 -2184
rect 774 -2218 808 -2184
rect 1008 -2218 1042 -2184
rect 1076 -2218 1110 -2184
rect 1144 -2218 1178 -2184
rect 1212 -2218 1246 -2184
rect 570 -2286 604 -2252
rect 1212 -2286 1246 -2252
rect 570 -2354 604 -2320
rect 570 -2422 604 -2388
rect 570 -2656 604 -2622
rect 570 -2724 604 -2690
rect 1212 -2354 1246 -2320
rect 1212 -2422 1246 -2388
rect 1212 -2656 1246 -2622
rect 1212 -2724 1246 -2690
rect 570 -2792 604 -2758
rect 1212 -2792 1246 -2758
rect 570 -2860 604 -2826
rect 638 -2860 672 -2826
rect 706 -2860 740 -2826
rect 774 -2860 808 -2826
rect 1008 -2860 1042 -2826
rect 1076 -2860 1110 -2826
rect 1144 -2860 1178 -2826
rect 1212 -2860 1246 -2826
rect 1390 -2218 1424 -2184
rect 1458 -2218 1492 -2184
rect 1526 -2218 1560 -2184
rect 1594 -2218 1628 -2184
rect 1828 -2218 1862 -2184
rect 1896 -2218 1930 -2184
rect 1964 -2218 1998 -2184
rect 2032 -2218 2066 -2184
rect 1390 -2286 1424 -2252
rect 2032 -2286 2066 -2252
rect 1390 -2354 1424 -2320
rect 1390 -2422 1424 -2388
rect 1390 -2656 1424 -2622
rect 1390 -2724 1424 -2690
rect 2032 -2354 2066 -2320
rect 2032 -2422 2066 -2388
rect 2032 -2656 2066 -2622
rect 2032 -2724 2066 -2690
rect 1390 -2792 1424 -2758
rect 2032 -2792 2066 -2758
rect 1390 -2860 1424 -2826
rect 1458 -2860 1492 -2826
rect 1526 -2860 1560 -2826
rect 1594 -2860 1628 -2826
rect 1828 -2860 1862 -2826
rect 1896 -2860 1930 -2826
rect 1964 -2860 1998 -2826
rect 2032 -2860 2066 -2826
rect 2210 -2218 2244 -2184
rect 2278 -2218 2312 -2184
rect 2346 -2218 2380 -2184
rect 2414 -2218 2448 -2184
rect 2648 -2218 2682 -2184
rect 2716 -2218 2750 -2184
rect 2784 -2218 2818 -2184
rect 2852 -2218 2886 -2184
rect 2210 -2286 2244 -2252
rect 2852 -2286 2886 -2252
rect 2210 -2354 2244 -2320
rect 2210 -2422 2244 -2388
rect 2210 -2656 2244 -2622
rect 2210 -2724 2244 -2690
rect 2852 -2354 2886 -2320
rect 2852 -2422 2886 -2388
rect 2852 -2656 2886 -2622
rect 2852 -2724 2886 -2690
rect 2210 -2792 2244 -2758
rect 2852 -2792 2886 -2758
rect 2210 -2860 2244 -2826
rect 2278 -2860 2312 -2826
rect 2346 -2860 2380 -2826
rect 2414 -2860 2448 -2826
rect 2648 -2860 2682 -2826
rect 2716 -2860 2750 -2826
rect 2784 -2860 2818 -2826
rect 2852 -2860 2886 -2826
rect 3030 -2218 3064 -2184
rect 3098 -2218 3132 -2184
rect 3166 -2218 3200 -2184
rect 3234 -2218 3268 -2184
rect 3468 -2218 3502 -2184
rect 3536 -2218 3570 -2184
rect 3604 -2218 3638 -2184
rect 3672 -2218 3706 -2184
rect 3030 -2286 3064 -2252
rect 3672 -2286 3706 -2252
rect 3030 -2354 3064 -2320
rect 3030 -2422 3064 -2388
rect 3030 -2656 3064 -2622
rect 3030 -2724 3064 -2690
rect 3672 -2354 3706 -2320
rect 3672 -2422 3706 -2388
rect 3672 -2656 3706 -2622
rect 3672 -2724 3706 -2690
rect 3030 -2792 3064 -2758
rect 3672 -2792 3706 -2758
rect 3030 -2860 3064 -2826
rect 3098 -2860 3132 -2826
rect 3166 -2860 3200 -2826
rect 3234 -2860 3268 -2826
rect 3468 -2860 3502 -2826
rect 3536 -2860 3570 -2826
rect 3604 -2860 3638 -2826
rect 3672 -2860 3706 -2826
rect 3850 -2218 3884 -2184
rect 3918 -2218 3952 -2184
rect 3986 -2218 4020 -2184
rect 4054 -2218 4088 -2184
rect 4288 -2218 4322 -2184
rect 4356 -2218 4390 -2184
rect 4424 -2218 4458 -2184
rect 4492 -2218 4526 -2184
rect 3850 -2286 3884 -2252
rect 4492 -2286 4526 -2252
rect 3850 -2354 3884 -2320
rect 3850 -2422 3884 -2388
rect 3850 -2656 3884 -2622
rect 3850 -2724 3884 -2690
rect 4492 -2354 4526 -2320
rect 4492 -2422 4526 -2388
rect 4492 -2656 4526 -2622
rect 4492 -2724 4526 -2690
rect 3850 -2792 3884 -2758
rect 4492 -2792 4526 -2758
rect 3850 -2860 3884 -2826
rect 3918 -2860 3952 -2826
rect 3986 -2860 4020 -2826
rect 4054 -2860 4088 -2826
rect 4288 -2860 4322 -2826
rect 4356 -2860 4390 -2826
rect 4424 -2860 4458 -2826
rect 4492 -2860 4526 -2826
rect 4670 -2218 4704 -2184
rect 4738 -2218 4772 -2184
rect 4806 -2218 4840 -2184
rect 4874 -2218 4908 -2184
rect 5108 -2218 5142 -2184
rect 5176 -2218 5210 -2184
rect 5244 -2218 5278 -2184
rect 5312 -2218 5346 -2184
rect 4670 -2286 4704 -2252
rect 5312 -2286 5346 -2252
rect 4670 -2354 4704 -2320
rect 4670 -2422 4704 -2388
rect 4670 -2656 4704 -2622
rect 4670 -2724 4704 -2690
rect 5312 -2354 5346 -2320
rect 5312 -2422 5346 -2388
rect 5312 -2656 5346 -2622
rect 5312 -2724 5346 -2690
rect 4670 -2792 4704 -2758
rect 5312 -2792 5346 -2758
rect 4670 -2860 4704 -2826
rect 4738 -2860 4772 -2826
rect 4806 -2860 4840 -2826
rect 4874 -2860 4908 -2826
rect 5108 -2860 5142 -2826
rect 5176 -2860 5210 -2826
rect 5244 -2860 5278 -2826
rect 5312 -2860 5346 -2826
rect 5490 -2218 5524 -2184
rect 5558 -2218 5592 -2184
rect 5626 -2218 5660 -2184
rect 5694 -2218 5728 -2184
rect 5928 -2218 5962 -2184
rect 5996 -2218 6030 -2184
rect 6064 -2218 6098 -2184
rect 6132 -2218 6166 -2184
rect 5490 -2286 5524 -2252
rect 6132 -2286 6166 -2252
rect 5490 -2354 5524 -2320
rect 5490 -2422 5524 -2388
rect 5490 -2656 5524 -2622
rect 5490 -2724 5524 -2690
rect 6132 -2354 6166 -2320
rect 6132 -2422 6166 -2388
rect 6132 -2656 6166 -2622
rect 6132 -2724 6166 -2690
rect 5490 -2792 5524 -2758
rect 6132 -2792 6166 -2758
rect 5490 -2860 5524 -2826
rect 5558 -2860 5592 -2826
rect 5626 -2860 5660 -2826
rect 5694 -2860 5728 -2826
rect 5928 -2860 5962 -2826
rect 5996 -2860 6030 -2826
rect 6064 -2860 6098 -2826
rect 6132 -2860 6166 -2826
rect 6310 -2218 6344 -2184
rect 6378 -2218 6412 -2184
rect 6446 -2218 6480 -2184
rect 6514 -2218 6548 -2184
rect 6748 -2218 6782 -2184
rect 6816 -2218 6850 -2184
rect 6884 -2218 6918 -2184
rect 6952 -2218 6986 -2184
rect 6310 -2286 6344 -2252
rect 6952 -2286 6986 -2252
rect 6310 -2354 6344 -2320
rect 6310 -2422 6344 -2388
rect 6310 -2656 6344 -2622
rect 6310 -2724 6344 -2690
rect 6952 -2354 6986 -2320
rect 6952 -2422 6986 -2388
rect 6952 -2656 6986 -2622
rect 6952 -2724 6986 -2690
rect 6310 -2792 6344 -2758
rect 6952 -2792 6986 -2758
rect 6310 -2860 6344 -2826
rect 6378 -2860 6412 -2826
rect 6446 -2860 6480 -2826
rect 6514 -2860 6548 -2826
rect 6748 -2860 6782 -2826
rect 6816 -2860 6850 -2826
rect 6884 -2860 6918 -2826
rect 6952 -2860 6986 -2826
rect -1070 -3038 -1036 -3004
rect -1002 -3038 -968 -3004
rect -934 -3038 -900 -3004
rect -866 -3038 -832 -3004
rect -632 -3038 -598 -3004
rect -564 -3038 -530 -3004
rect -496 -3038 -462 -3004
rect -428 -3038 -394 -3004
rect -1070 -3106 -1036 -3072
rect -428 -3106 -394 -3072
rect -1070 -3174 -1036 -3140
rect -1070 -3242 -1036 -3208
rect -1070 -3476 -1036 -3442
rect -1070 -3544 -1036 -3510
rect -428 -3174 -394 -3140
rect -428 -3242 -394 -3208
rect -428 -3476 -394 -3442
rect -428 -3544 -394 -3510
rect -1070 -3612 -1036 -3578
rect -428 -3612 -394 -3578
rect -1070 -3680 -1036 -3646
rect -1002 -3680 -968 -3646
rect -934 -3680 -900 -3646
rect -866 -3680 -832 -3646
rect -632 -3680 -598 -3646
rect -564 -3680 -530 -3646
rect -496 -3680 -462 -3646
rect -428 -3680 -394 -3646
rect -250 -3038 -216 -3004
rect -182 -3038 -148 -3004
rect -114 -3038 -80 -3004
rect -46 -3038 -12 -3004
rect 188 -3038 222 -3004
rect 256 -3038 290 -3004
rect 324 -3038 358 -3004
rect 392 -3038 426 -3004
rect -250 -3106 -216 -3072
rect 392 -3106 426 -3072
rect -250 -3174 -216 -3140
rect -250 -3242 -216 -3208
rect -250 -3476 -216 -3442
rect -250 -3544 -216 -3510
rect 392 -3174 426 -3140
rect 392 -3242 426 -3208
rect 392 -3476 426 -3442
rect 392 -3544 426 -3510
rect -250 -3612 -216 -3578
rect 392 -3612 426 -3578
rect -250 -3680 -216 -3646
rect -182 -3680 -148 -3646
rect -114 -3680 -80 -3646
rect -46 -3680 -12 -3646
rect 188 -3680 222 -3646
rect 256 -3680 290 -3646
rect 324 -3680 358 -3646
rect 392 -3680 426 -3646
rect 570 -3038 604 -3004
rect 638 -3038 672 -3004
rect 706 -3038 740 -3004
rect 774 -3038 808 -3004
rect 1008 -3038 1042 -3004
rect 1076 -3038 1110 -3004
rect 1144 -3038 1178 -3004
rect 1212 -3038 1246 -3004
rect 570 -3106 604 -3072
rect 1212 -3106 1246 -3072
rect 570 -3174 604 -3140
rect 570 -3242 604 -3208
rect 570 -3476 604 -3442
rect 570 -3544 604 -3510
rect 1212 -3174 1246 -3140
rect 1212 -3242 1246 -3208
rect 1212 -3476 1246 -3442
rect 1212 -3544 1246 -3510
rect 570 -3612 604 -3578
rect 1212 -3612 1246 -3578
rect 570 -3680 604 -3646
rect 638 -3680 672 -3646
rect 706 -3680 740 -3646
rect 774 -3680 808 -3646
rect 1008 -3680 1042 -3646
rect 1076 -3680 1110 -3646
rect 1144 -3680 1178 -3646
rect 1212 -3680 1246 -3646
rect 1390 -3038 1424 -3004
rect 1458 -3038 1492 -3004
rect 1526 -3038 1560 -3004
rect 1594 -3038 1628 -3004
rect 1828 -3038 1862 -3004
rect 1896 -3038 1930 -3004
rect 1964 -3038 1998 -3004
rect 2032 -3038 2066 -3004
rect 1390 -3106 1424 -3072
rect 2032 -3106 2066 -3072
rect 1390 -3174 1424 -3140
rect 1390 -3242 1424 -3208
rect 1390 -3476 1424 -3442
rect 1390 -3544 1424 -3510
rect 2032 -3174 2066 -3140
rect 2032 -3242 2066 -3208
rect 2032 -3476 2066 -3442
rect 2032 -3544 2066 -3510
rect 1390 -3612 1424 -3578
rect 2032 -3612 2066 -3578
rect 1390 -3680 1424 -3646
rect 1458 -3680 1492 -3646
rect 1526 -3680 1560 -3646
rect 1594 -3680 1628 -3646
rect 1828 -3680 1862 -3646
rect 1896 -3680 1930 -3646
rect 1964 -3680 1998 -3646
rect 2032 -3680 2066 -3646
rect 2210 -3038 2244 -3004
rect 2278 -3038 2312 -3004
rect 2346 -3038 2380 -3004
rect 2414 -3038 2448 -3004
rect 2648 -3038 2682 -3004
rect 2716 -3038 2750 -3004
rect 2784 -3038 2818 -3004
rect 2852 -3038 2886 -3004
rect 2210 -3106 2244 -3072
rect 2852 -3106 2886 -3072
rect 2210 -3174 2244 -3140
rect 2210 -3242 2244 -3208
rect 2210 -3476 2244 -3442
rect 2210 -3544 2244 -3510
rect 2852 -3174 2886 -3140
rect 2852 -3242 2886 -3208
rect 2852 -3476 2886 -3442
rect 2852 -3544 2886 -3510
rect 2210 -3612 2244 -3578
rect 2852 -3612 2886 -3578
rect 2210 -3680 2244 -3646
rect 2278 -3680 2312 -3646
rect 2346 -3680 2380 -3646
rect 2414 -3680 2448 -3646
rect 2648 -3680 2682 -3646
rect 2716 -3680 2750 -3646
rect 2784 -3680 2818 -3646
rect 2852 -3680 2886 -3646
rect 3030 -3038 3064 -3004
rect 3098 -3038 3132 -3004
rect 3166 -3038 3200 -3004
rect 3234 -3038 3268 -3004
rect 3468 -3038 3502 -3004
rect 3536 -3038 3570 -3004
rect 3604 -3038 3638 -3004
rect 3672 -3038 3706 -3004
rect 3030 -3106 3064 -3072
rect 3672 -3106 3706 -3072
rect 3030 -3174 3064 -3140
rect 3030 -3242 3064 -3208
rect 3030 -3476 3064 -3442
rect 3030 -3544 3064 -3510
rect 3672 -3174 3706 -3140
rect 3672 -3242 3706 -3208
rect 3672 -3476 3706 -3442
rect 3672 -3544 3706 -3510
rect 3030 -3612 3064 -3578
rect 3672 -3612 3706 -3578
rect 3030 -3680 3064 -3646
rect 3098 -3680 3132 -3646
rect 3166 -3680 3200 -3646
rect 3234 -3680 3268 -3646
rect 3468 -3680 3502 -3646
rect 3536 -3680 3570 -3646
rect 3604 -3680 3638 -3646
rect 3672 -3680 3706 -3646
rect 3850 -3038 3884 -3004
rect 3918 -3038 3952 -3004
rect 3986 -3038 4020 -3004
rect 4054 -3038 4088 -3004
rect 4288 -3038 4322 -3004
rect 4356 -3038 4390 -3004
rect 4424 -3038 4458 -3004
rect 4492 -3038 4526 -3004
rect 3850 -3106 3884 -3072
rect 4492 -3106 4526 -3072
rect 3850 -3174 3884 -3140
rect 3850 -3242 3884 -3208
rect 3850 -3476 3884 -3442
rect 3850 -3544 3884 -3510
rect 4492 -3174 4526 -3140
rect 4492 -3242 4526 -3208
rect 4492 -3476 4526 -3442
rect 4492 -3544 4526 -3510
rect 3850 -3612 3884 -3578
rect 4492 -3612 4526 -3578
rect 3850 -3680 3884 -3646
rect 3918 -3680 3952 -3646
rect 3986 -3680 4020 -3646
rect 4054 -3680 4088 -3646
rect 4288 -3680 4322 -3646
rect 4356 -3680 4390 -3646
rect 4424 -3680 4458 -3646
rect 4492 -3680 4526 -3646
rect 4670 -3038 4704 -3004
rect 4738 -3038 4772 -3004
rect 4806 -3038 4840 -3004
rect 4874 -3038 4908 -3004
rect 5108 -3038 5142 -3004
rect 5176 -3038 5210 -3004
rect 5244 -3038 5278 -3004
rect 5312 -3038 5346 -3004
rect 4670 -3106 4704 -3072
rect 5312 -3106 5346 -3072
rect 4670 -3174 4704 -3140
rect 4670 -3242 4704 -3208
rect 4670 -3476 4704 -3442
rect 4670 -3544 4704 -3510
rect 5312 -3174 5346 -3140
rect 5312 -3242 5346 -3208
rect 5312 -3476 5346 -3442
rect 5312 -3544 5346 -3510
rect 4670 -3612 4704 -3578
rect 5312 -3612 5346 -3578
rect 4670 -3680 4704 -3646
rect 4738 -3680 4772 -3646
rect 4806 -3680 4840 -3646
rect 4874 -3680 4908 -3646
rect 5108 -3680 5142 -3646
rect 5176 -3680 5210 -3646
rect 5244 -3680 5278 -3646
rect 5312 -3680 5346 -3646
rect 5490 -3038 5524 -3004
rect 5558 -3038 5592 -3004
rect 5626 -3038 5660 -3004
rect 5694 -3038 5728 -3004
rect 5928 -3038 5962 -3004
rect 5996 -3038 6030 -3004
rect 6064 -3038 6098 -3004
rect 6132 -3038 6166 -3004
rect 5490 -3106 5524 -3072
rect 6132 -3106 6166 -3072
rect 5490 -3174 5524 -3140
rect 5490 -3242 5524 -3208
rect 5490 -3476 5524 -3442
rect 5490 -3544 5524 -3510
rect 6132 -3174 6166 -3140
rect 6132 -3242 6166 -3208
rect 6132 -3476 6166 -3442
rect 6132 -3544 6166 -3510
rect 5490 -3612 5524 -3578
rect 6132 -3612 6166 -3578
rect 5490 -3680 5524 -3646
rect 5558 -3680 5592 -3646
rect 5626 -3680 5660 -3646
rect 5694 -3680 5728 -3646
rect 5928 -3680 5962 -3646
rect 5996 -3680 6030 -3646
rect 6064 -3680 6098 -3646
rect 6132 -3680 6166 -3646
rect 6310 -3038 6344 -3004
rect 6378 -3038 6412 -3004
rect 6446 -3038 6480 -3004
rect 6514 -3038 6548 -3004
rect 6748 -3038 6782 -3004
rect 6816 -3038 6850 -3004
rect 6884 -3038 6918 -3004
rect 6952 -3038 6986 -3004
rect 6310 -3106 6344 -3072
rect 6952 -3106 6986 -3072
rect 6310 -3174 6344 -3140
rect 6310 -3242 6344 -3208
rect 6310 -3476 6344 -3442
rect 6310 -3544 6344 -3510
rect 6952 -3174 6986 -3140
rect 6952 -3242 6986 -3208
rect 6952 -3476 6986 -3442
rect 6952 -3544 6986 -3510
rect 6310 -3612 6344 -3578
rect 6952 -3612 6986 -3578
rect 6310 -3680 6344 -3646
rect 6378 -3680 6412 -3646
rect 6446 -3680 6480 -3646
rect 6514 -3680 6548 -3646
rect 6748 -3680 6782 -3646
rect 6816 -3680 6850 -3646
rect 6884 -3680 6918 -3646
rect 6952 -3680 6986 -3646
rect -1070 -3858 -1036 -3824
rect -1002 -3858 -968 -3824
rect -934 -3858 -900 -3824
rect -866 -3858 -832 -3824
rect -632 -3858 -598 -3824
rect -564 -3858 -530 -3824
rect -496 -3858 -462 -3824
rect -428 -3858 -394 -3824
rect -1070 -3926 -1036 -3892
rect -428 -3926 -394 -3892
rect -1070 -3994 -1036 -3960
rect -1070 -4062 -1036 -4028
rect -1070 -4296 -1036 -4262
rect -1070 -4364 -1036 -4330
rect -428 -3994 -394 -3960
rect -428 -4062 -394 -4028
rect -428 -4296 -394 -4262
rect -428 -4364 -394 -4330
rect -1070 -4432 -1036 -4398
rect -428 -4432 -394 -4398
rect -1070 -4500 -1036 -4466
rect -1002 -4500 -968 -4466
rect -934 -4500 -900 -4466
rect -866 -4500 -832 -4466
rect -632 -4500 -598 -4466
rect -564 -4500 -530 -4466
rect -496 -4500 -462 -4466
rect -428 -4500 -394 -4466
rect -250 -3858 -216 -3824
rect -182 -3858 -148 -3824
rect -114 -3858 -80 -3824
rect -46 -3858 -12 -3824
rect 188 -3858 222 -3824
rect 256 -3858 290 -3824
rect 324 -3858 358 -3824
rect 392 -3858 426 -3824
rect -250 -3926 -216 -3892
rect 392 -3926 426 -3892
rect -250 -3994 -216 -3960
rect -250 -4062 -216 -4028
rect -250 -4296 -216 -4262
rect -250 -4364 -216 -4330
rect 392 -3994 426 -3960
rect 392 -4062 426 -4028
rect 392 -4296 426 -4262
rect 392 -4364 426 -4330
rect -250 -4432 -216 -4398
rect 392 -4432 426 -4398
rect -250 -4500 -216 -4466
rect -182 -4500 -148 -4466
rect -114 -4500 -80 -4466
rect -46 -4500 -12 -4466
rect 188 -4500 222 -4466
rect 256 -4500 290 -4466
rect 324 -4500 358 -4466
rect 392 -4500 426 -4466
rect 570 -3858 604 -3824
rect 638 -3858 672 -3824
rect 706 -3858 740 -3824
rect 774 -3858 808 -3824
rect 1008 -3858 1042 -3824
rect 1076 -3858 1110 -3824
rect 1144 -3858 1178 -3824
rect 1212 -3858 1246 -3824
rect 570 -3926 604 -3892
rect 1212 -3926 1246 -3892
rect 570 -3994 604 -3960
rect 570 -4062 604 -4028
rect 570 -4296 604 -4262
rect 570 -4364 604 -4330
rect 1212 -3994 1246 -3960
rect 1212 -4062 1246 -4028
rect 1212 -4296 1246 -4262
rect 1212 -4364 1246 -4330
rect 570 -4432 604 -4398
rect 1212 -4432 1246 -4398
rect 570 -4500 604 -4466
rect 638 -4500 672 -4466
rect 706 -4500 740 -4466
rect 774 -4500 808 -4466
rect 1008 -4500 1042 -4466
rect 1076 -4500 1110 -4466
rect 1144 -4500 1178 -4466
rect 1212 -4500 1246 -4466
rect 1390 -3858 1424 -3824
rect 1458 -3858 1492 -3824
rect 1526 -3858 1560 -3824
rect 1594 -3858 1628 -3824
rect 1828 -3858 1862 -3824
rect 1896 -3858 1930 -3824
rect 1964 -3858 1998 -3824
rect 2032 -3858 2066 -3824
rect 1390 -3926 1424 -3892
rect 2032 -3926 2066 -3892
rect 1390 -3994 1424 -3960
rect 1390 -4062 1424 -4028
rect 1390 -4296 1424 -4262
rect 1390 -4364 1424 -4330
rect 2032 -3994 2066 -3960
rect 2032 -4062 2066 -4028
rect 2032 -4296 2066 -4262
rect 2032 -4364 2066 -4330
rect 1390 -4432 1424 -4398
rect 2032 -4432 2066 -4398
rect 1390 -4500 1424 -4466
rect 1458 -4500 1492 -4466
rect 1526 -4500 1560 -4466
rect 1594 -4500 1628 -4466
rect 1828 -4500 1862 -4466
rect 1896 -4500 1930 -4466
rect 1964 -4500 1998 -4466
rect 2032 -4500 2066 -4466
rect 2210 -3858 2244 -3824
rect 2278 -3858 2312 -3824
rect 2346 -3858 2380 -3824
rect 2414 -3858 2448 -3824
rect 2648 -3858 2682 -3824
rect 2716 -3858 2750 -3824
rect 2784 -3858 2818 -3824
rect 2852 -3858 2886 -3824
rect 2210 -3926 2244 -3892
rect 2852 -3926 2886 -3892
rect 2210 -3994 2244 -3960
rect 2210 -4062 2244 -4028
rect 2210 -4296 2244 -4262
rect 2210 -4364 2244 -4330
rect 2852 -3994 2886 -3960
rect 2852 -4062 2886 -4028
rect 2852 -4296 2886 -4262
rect 2852 -4364 2886 -4330
rect 2210 -4432 2244 -4398
rect 2852 -4432 2886 -4398
rect 2210 -4500 2244 -4466
rect 2278 -4500 2312 -4466
rect 2346 -4500 2380 -4466
rect 2414 -4500 2448 -4466
rect 2648 -4500 2682 -4466
rect 2716 -4500 2750 -4466
rect 2784 -4500 2818 -4466
rect 2852 -4500 2886 -4466
rect 3030 -3858 3064 -3824
rect 3098 -3858 3132 -3824
rect 3166 -3858 3200 -3824
rect 3234 -3858 3268 -3824
rect 3468 -3858 3502 -3824
rect 3536 -3858 3570 -3824
rect 3604 -3858 3638 -3824
rect 3672 -3858 3706 -3824
rect 3030 -3926 3064 -3892
rect 3672 -3926 3706 -3892
rect 3030 -3994 3064 -3960
rect 3030 -4062 3064 -4028
rect 3030 -4296 3064 -4262
rect 3030 -4364 3064 -4330
rect 3672 -3994 3706 -3960
rect 3672 -4062 3706 -4028
rect 3672 -4296 3706 -4262
rect 3672 -4364 3706 -4330
rect 3030 -4432 3064 -4398
rect 3672 -4432 3706 -4398
rect 3030 -4500 3064 -4466
rect 3098 -4500 3132 -4466
rect 3166 -4500 3200 -4466
rect 3234 -4500 3268 -4466
rect 3468 -4500 3502 -4466
rect 3536 -4500 3570 -4466
rect 3604 -4500 3638 -4466
rect 3672 -4500 3706 -4466
rect 3850 -3858 3884 -3824
rect 3918 -3858 3952 -3824
rect 3986 -3858 4020 -3824
rect 4054 -3858 4088 -3824
rect 4288 -3858 4322 -3824
rect 4356 -3858 4390 -3824
rect 4424 -3858 4458 -3824
rect 4492 -3858 4526 -3824
rect 3850 -3926 3884 -3892
rect 4492 -3926 4526 -3892
rect 3850 -3994 3884 -3960
rect 3850 -4062 3884 -4028
rect 3850 -4296 3884 -4262
rect 3850 -4364 3884 -4330
rect 4492 -3994 4526 -3960
rect 4492 -4062 4526 -4028
rect 4492 -4296 4526 -4262
rect 4492 -4364 4526 -4330
rect 3850 -4432 3884 -4398
rect 4492 -4432 4526 -4398
rect 3850 -4500 3884 -4466
rect 3918 -4500 3952 -4466
rect 3986 -4500 4020 -4466
rect 4054 -4500 4088 -4466
rect 4288 -4500 4322 -4466
rect 4356 -4500 4390 -4466
rect 4424 -4500 4458 -4466
rect 4492 -4500 4526 -4466
rect 4670 -3858 4704 -3824
rect 4738 -3858 4772 -3824
rect 4806 -3858 4840 -3824
rect 4874 -3858 4908 -3824
rect 5108 -3858 5142 -3824
rect 5176 -3858 5210 -3824
rect 5244 -3858 5278 -3824
rect 5312 -3858 5346 -3824
rect 4670 -3926 4704 -3892
rect 5312 -3926 5346 -3892
rect 4670 -3994 4704 -3960
rect 4670 -4062 4704 -4028
rect 4670 -4296 4704 -4262
rect 4670 -4364 4704 -4330
rect 5312 -3994 5346 -3960
rect 5312 -4062 5346 -4028
rect 5312 -4296 5346 -4262
rect 5312 -4364 5346 -4330
rect 4670 -4432 4704 -4398
rect 5312 -4432 5346 -4398
rect 4670 -4500 4704 -4466
rect 4738 -4500 4772 -4466
rect 4806 -4500 4840 -4466
rect 4874 -4500 4908 -4466
rect 5108 -4500 5142 -4466
rect 5176 -4500 5210 -4466
rect 5244 -4500 5278 -4466
rect 5312 -4500 5346 -4466
rect 5490 -3858 5524 -3824
rect 5558 -3858 5592 -3824
rect 5626 -3858 5660 -3824
rect 5694 -3858 5728 -3824
rect 5928 -3858 5962 -3824
rect 5996 -3858 6030 -3824
rect 6064 -3858 6098 -3824
rect 6132 -3858 6166 -3824
rect 5490 -3926 5524 -3892
rect 6132 -3926 6166 -3892
rect 5490 -3994 5524 -3960
rect 5490 -4062 5524 -4028
rect 5490 -4296 5524 -4262
rect 5490 -4364 5524 -4330
rect 6132 -3994 6166 -3960
rect 6132 -4062 6166 -4028
rect 6132 -4296 6166 -4262
rect 6132 -4364 6166 -4330
rect 5490 -4432 5524 -4398
rect 6132 -4432 6166 -4398
rect 5490 -4500 5524 -4466
rect 5558 -4500 5592 -4466
rect 5626 -4500 5660 -4466
rect 5694 -4500 5728 -4466
rect 5928 -4500 5962 -4466
rect 5996 -4500 6030 -4466
rect 6064 -4500 6098 -4466
rect 6132 -4500 6166 -4466
rect 6310 -3858 6344 -3824
rect 6378 -3858 6412 -3824
rect 6446 -3858 6480 -3824
rect 6514 -3858 6548 -3824
rect 6748 -3858 6782 -3824
rect 6816 -3858 6850 -3824
rect 6884 -3858 6918 -3824
rect 6952 -3858 6986 -3824
rect 6310 -3926 6344 -3892
rect 6952 -3926 6986 -3892
rect 6310 -3994 6344 -3960
rect 6310 -4062 6344 -4028
rect 6310 -4296 6344 -4262
rect 6310 -4364 6344 -4330
rect 6952 -3994 6986 -3960
rect 6952 -4062 6986 -4028
rect 6952 -4296 6986 -4262
rect 6952 -4364 6986 -4330
rect 6310 -4432 6344 -4398
rect 6952 -4432 6986 -4398
rect 6310 -4500 6344 -4466
rect 6378 -4500 6412 -4466
rect 6446 -4500 6480 -4466
rect 6514 -4500 6548 -4466
rect 6748 -4500 6782 -4466
rect 6816 -4500 6850 -4466
rect 6884 -4500 6918 -4466
rect 6952 -4500 6986 -4466
<< nsubdiffcont >>
rect 7660 4300 7700 6240
rect 7660 2090 7700 4030
rect -917 -731 -883 -697
rect -849 -731 -815 -697
rect -649 -731 -615 -697
rect -581 -731 -547 -697
rect -917 -799 -883 -765
rect -581 -799 -547 -765
rect -917 -999 -883 -965
rect -581 -999 -547 -965
rect -917 -1067 -883 -1033
rect -849 -1067 -815 -1033
rect -649 -1067 -615 -1033
rect -581 -1067 -547 -1033
rect -97 -731 -63 -697
rect -29 -731 5 -697
rect 171 -731 205 -697
rect 239 -731 273 -697
rect -97 -799 -63 -765
rect 239 -799 273 -765
rect -97 -999 -63 -965
rect 239 -999 273 -965
rect -97 -1067 -63 -1033
rect -29 -1067 5 -1033
rect 171 -1067 205 -1033
rect 239 -1067 273 -1033
rect 723 -731 757 -697
rect 791 -731 825 -697
rect 991 -731 1025 -697
rect 1059 -731 1093 -697
rect 723 -799 757 -765
rect 1059 -799 1093 -765
rect 723 -999 757 -965
rect 1059 -999 1093 -965
rect 723 -1067 757 -1033
rect 791 -1067 825 -1033
rect 991 -1067 1025 -1033
rect 1059 -1067 1093 -1033
rect 1543 -731 1577 -697
rect 1611 -731 1645 -697
rect 1811 -731 1845 -697
rect 1879 -731 1913 -697
rect 1543 -799 1577 -765
rect 1879 -799 1913 -765
rect 1543 -999 1577 -965
rect 1879 -999 1913 -965
rect 1543 -1067 1577 -1033
rect 1611 -1067 1645 -1033
rect 1811 -1067 1845 -1033
rect 1879 -1067 1913 -1033
rect 2363 -731 2397 -697
rect 2431 -731 2465 -697
rect 2631 -731 2665 -697
rect 2699 -731 2733 -697
rect 2363 -799 2397 -765
rect 2699 -799 2733 -765
rect 2363 -999 2397 -965
rect 2699 -999 2733 -965
rect 2363 -1067 2397 -1033
rect 2431 -1067 2465 -1033
rect 2631 -1067 2665 -1033
rect 2699 -1067 2733 -1033
rect 3183 -731 3217 -697
rect 3251 -731 3285 -697
rect 3451 -731 3485 -697
rect 3519 -731 3553 -697
rect 3183 -799 3217 -765
rect 3519 -799 3553 -765
rect 3183 -999 3217 -965
rect 3519 -999 3553 -965
rect 3183 -1067 3217 -1033
rect 3251 -1067 3285 -1033
rect 3451 -1067 3485 -1033
rect 3519 -1067 3553 -1033
rect 4003 -731 4037 -697
rect 4071 -731 4105 -697
rect 4271 -731 4305 -697
rect 4339 -731 4373 -697
rect 4003 -799 4037 -765
rect 4339 -799 4373 -765
rect 4003 -999 4037 -965
rect 4339 -999 4373 -965
rect 4003 -1067 4037 -1033
rect 4071 -1067 4105 -1033
rect 4271 -1067 4305 -1033
rect 4339 -1067 4373 -1033
rect 4823 -731 4857 -697
rect 4891 -731 4925 -697
rect 5091 -731 5125 -697
rect 5159 -731 5193 -697
rect 4823 -799 4857 -765
rect 5159 -799 5193 -765
rect 4823 -999 4857 -965
rect 5159 -999 5193 -965
rect 4823 -1067 4857 -1033
rect 4891 -1067 4925 -1033
rect 5091 -1067 5125 -1033
rect 5159 -1067 5193 -1033
rect 5643 -731 5677 -697
rect 5711 -731 5745 -697
rect 5911 -731 5945 -697
rect 5979 -731 6013 -697
rect 5643 -799 5677 -765
rect 5979 -799 6013 -765
rect 5643 -999 5677 -965
rect 5979 -999 6013 -965
rect 5643 -1067 5677 -1033
rect 5711 -1067 5745 -1033
rect 5911 -1067 5945 -1033
rect 5979 -1067 6013 -1033
rect 6463 -731 6497 -697
rect 6531 -731 6565 -697
rect 6731 -731 6765 -697
rect 6799 -731 6833 -697
rect 6463 -799 6497 -765
rect 6799 -799 6833 -765
rect 6463 -999 6497 -965
rect 6799 -999 6833 -965
rect 6463 -1067 6497 -1033
rect 6531 -1067 6565 -1033
rect 6731 -1067 6765 -1033
rect 6799 -1067 6833 -1033
rect 7313 -731 7347 -697
rect 7381 -731 7415 -697
rect 7581 -731 7615 -697
rect 7649 -731 7683 -697
rect 7313 -799 7347 -765
rect 7649 -799 7683 -765
rect 7313 -999 7347 -965
rect 7649 -999 7683 -965
rect 7313 -1067 7347 -1033
rect 7381 -1067 7415 -1033
rect 7581 -1067 7615 -1033
rect 7649 -1067 7683 -1033
rect -917 -1551 -883 -1517
rect -849 -1551 -815 -1517
rect -649 -1551 -615 -1517
rect -581 -1551 -547 -1517
rect -917 -1619 -883 -1585
rect -581 -1619 -547 -1585
rect -917 -1819 -883 -1785
rect -581 -1819 -547 -1785
rect -917 -1887 -883 -1853
rect -849 -1887 -815 -1853
rect -649 -1887 -615 -1853
rect -581 -1887 -547 -1853
rect -97 -1551 -63 -1517
rect -29 -1551 5 -1517
rect 171 -1551 205 -1517
rect 239 -1551 273 -1517
rect -97 -1619 -63 -1585
rect 239 -1619 273 -1585
rect -97 -1819 -63 -1785
rect 239 -1819 273 -1785
rect -97 -1887 -63 -1853
rect -29 -1887 5 -1853
rect 171 -1887 205 -1853
rect 239 -1887 273 -1853
rect 723 -1551 757 -1517
rect 791 -1551 825 -1517
rect 991 -1551 1025 -1517
rect 1059 -1551 1093 -1517
rect 723 -1619 757 -1585
rect 1059 -1619 1093 -1585
rect 723 -1819 757 -1785
rect 1059 -1819 1093 -1785
rect 723 -1887 757 -1853
rect 791 -1887 825 -1853
rect 991 -1887 1025 -1853
rect 1059 -1887 1093 -1853
rect 1543 -1551 1577 -1517
rect 1611 -1551 1645 -1517
rect 1811 -1551 1845 -1517
rect 1879 -1551 1913 -1517
rect 1543 -1619 1577 -1585
rect 1879 -1619 1913 -1585
rect 1543 -1819 1577 -1785
rect 1879 -1819 1913 -1785
rect 1543 -1887 1577 -1853
rect 1611 -1887 1645 -1853
rect 1811 -1887 1845 -1853
rect 1879 -1887 1913 -1853
rect 2363 -1551 2397 -1517
rect 2431 -1551 2465 -1517
rect 2631 -1551 2665 -1517
rect 2699 -1551 2733 -1517
rect 2363 -1619 2397 -1585
rect 2699 -1619 2733 -1585
rect 2363 -1819 2397 -1785
rect 2699 -1819 2733 -1785
rect 2363 -1887 2397 -1853
rect 2431 -1887 2465 -1853
rect 2631 -1887 2665 -1853
rect 2699 -1887 2733 -1853
rect 3183 -1551 3217 -1517
rect 3251 -1551 3285 -1517
rect 3451 -1551 3485 -1517
rect 3519 -1551 3553 -1517
rect 3183 -1619 3217 -1585
rect 3519 -1619 3553 -1585
rect 3183 -1819 3217 -1785
rect 3519 -1819 3553 -1785
rect 3183 -1887 3217 -1853
rect 3251 -1887 3285 -1853
rect 3451 -1887 3485 -1853
rect 3519 -1887 3553 -1853
rect 4003 -1551 4037 -1517
rect 4071 -1551 4105 -1517
rect 4271 -1551 4305 -1517
rect 4339 -1551 4373 -1517
rect 4003 -1619 4037 -1585
rect 4339 -1619 4373 -1585
rect 4003 -1819 4037 -1785
rect 4339 -1819 4373 -1785
rect 4003 -1887 4037 -1853
rect 4071 -1887 4105 -1853
rect 4271 -1887 4305 -1853
rect 4339 -1887 4373 -1853
rect 4823 -1551 4857 -1517
rect 4891 -1551 4925 -1517
rect 5091 -1551 5125 -1517
rect 5159 -1551 5193 -1517
rect 4823 -1619 4857 -1585
rect 5159 -1619 5193 -1585
rect 4823 -1819 4857 -1785
rect 5159 -1819 5193 -1785
rect 4823 -1887 4857 -1853
rect 4891 -1887 4925 -1853
rect 5091 -1887 5125 -1853
rect 5159 -1887 5193 -1853
rect 5643 -1551 5677 -1517
rect 5711 -1551 5745 -1517
rect 5911 -1551 5945 -1517
rect 5979 -1551 6013 -1517
rect 5643 -1619 5677 -1585
rect 5979 -1619 6013 -1585
rect 5643 -1819 5677 -1785
rect 5979 -1819 6013 -1785
rect 5643 -1887 5677 -1853
rect 5711 -1887 5745 -1853
rect 5911 -1887 5945 -1853
rect 5979 -1887 6013 -1853
rect 6463 -1551 6497 -1517
rect 6531 -1551 6565 -1517
rect 6731 -1551 6765 -1517
rect 6799 -1551 6833 -1517
rect 6463 -1619 6497 -1585
rect 6799 -1619 6833 -1585
rect 6463 -1819 6497 -1785
rect 6799 -1819 6833 -1785
rect 6463 -1887 6497 -1853
rect 6531 -1887 6565 -1853
rect 6731 -1887 6765 -1853
rect 6799 -1887 6833 -1853
rect -917 -2371 -883 -2337
rect -849 -2371 -815 -2337
rect -649 -2371 -615 -2337
rect -581 -2371 -547 -2337
rect -917 -2439 -883 -2405
rect -581 -2439 -547 -2405
rect -917 -2639 -883 -2605
rect -581 -2639 -547 -2605
rect -917 -2707 -883 -2673
rect -849 -2707 -815 -2673
rect -649 -2707 -615 -2673
rect -581 -2707 -547 -2673
rect -97 -2371 -63 -2337
rect -29 -2371 5 -2337
rect 171 -2371 205 -2337
rect 239 -2371 273 -2337
rect -97 -2439 -63 -2405
rect 239 -2439 273 -2405
rect -97 -2639 -63 -2605
rect 239 -2639 273 -2605
rect -97 -2707 -63 -2673
rect -29 -2707 5 -2673
rect 171 -2707 205 -2673
rect 239 -2707 273 -2673
rect 723 -2371 757 -2337
rect 791 -2371 825 -2337
rect 991 -2371 1025 -2337
rect 1059 -2371 1093 -2337
rect 723 -2439 757 -2405
rect 1059 -2439 1093 -2405
rect 723 -2639 757 -2605
rect 1059 -2639 1093 -2605
rect 723 -2707 757 -2673
rect 791 -2707 825 -2673
rect 991 -2707 1025 -2673
rect 1059 -2707 1093 -2673
rect 1543 -2371 1577 -2337
rect 1611 -2371 1645 -2337
rect 1811 -2371 1845 -2337
rect 1879 -2371 1913 -2337
rect 1543 -2439 1577 -2405
rect 1879 -2439 1913 -2405
rect 1543 -2639 1577 -2605
rect 1879 -2639 1913 -2605
rect 1543 -2707 1577 -2673
rect 1611 -2707 1645 -2673
rect 1811 -2707 1845 -2673
rect 1879 -2707 1913 -2673
rect 2363 -2371 2397 -2337
rect 2431 -2371 2465 -2337
rect 2631 -2371 2665 -2337
rect 2699 -2371 2733 -2337
rect 2363 -2439 2397 -2405
rect 2699 -2439 2733 -2405
rect 2363 -2639 2397 -2605
rect 2699 -2639 2733 -2605
rect 2363 -2707 2397 -2673
rect 2431 -2707 2465 -2673
rect 2631 -2707 2665 -2673
rect 2699 -2707 2733 -2673
rect 3183 -2371 3217 -2337
rect 3251 -2371 3285 -2337
rect 3451 -2371 3485 -2337
rect 3519 -2371 3553 -2337
rect 3183 -2439 3217 -2405
rect 3519 -2439 3553 -2405
rect 3183 -2639 3217 -2605
rect 3519 -2639 3553 -2605
rect 3183 -2707 3217 -2673
rect 3251 -2707 3285 -2673
rect 3451 -2707 3485 -2673
rect 3519 -2707 3553 -2673
rect 4003 -2371 4037 -2337
rect 4071 -2371 4105 -2337
rect 4271 -2371 4305 -2337
rect 4339 -2371 4373 -2337
rect 4003 -2439 4037 -2405
rect 4339 -2439 4373 -2405
rect 4003 -2639 4037 -2605
rect 4339 -2639 4373 -2605
rect 4003 -2707 4037 -2673
rect 4071 -2707 4105 -2673
rect 4271 -2707 4305 -2673
rect 4339 -2707 4373 -2673
rect 4823 -2371 4857 -2337
rect 4891 -2371 4925 -2337
rect 5091 -2371 5125 -2337
rect 5159 -2371 5193 -2337
rect 4823 -2439 4857 -2405
rect 5159 -2439 5193 -2405
rect 4823 -2639 4857 -2605
rect 5159 -2639 5193 -2605
rect 4823 -2707 4857 -2673
rect 4891 -2707 4925 -2673
rect 5091 -2707 5125 -2673
rect 5159 -2707 5193 -2673
rect 5643 -2371 5677 -2337
rect 5711 -2371 5745 -2337
rect 5911 -2371 5945 -2337
rect 5979 -2371 6013 -2337
rect 5643 -2439 5677 -2405
rect 5979 -2439 6013 -2405
rect 5643 -2639 5677 -2605
rect 5979 -2639 6013 -2605
rect 5643 -2707 5677 -2673
rect 5711 -2707 5745 -2673
rect 5911 -2707 5945 -2673
rect 5979 -2707 6013 -2673
rect 6463 -2371 6497 -2337
rect 6531 -2371 6565 -2337
rect 6731 -2371 6765 -2337
rect 6799 -2371 6833 -2337
rect 6463 -2439 6497 -2405
rect 6799 -2439 6833 -2405
rect 6463 -2639 6497 -2605
rect 6799 -2639 6833 -2605
rect 6463 -2707 6497 -2673
rect 6531 -2707 6565 -2673
rect 6731 -2707 6765 -2673
rect 6799 -2707 6833 -2673
rect -917 -3191 -883 -3157
rect -849 -3191 -815 -3157
rect -649 -3191 -615 -3157
rect -581 -3191 -547 -3157
rect -917 -3259 -883 -3225
rect -581 -3259 -547 -3225
rect -917 -3459 -883 -3425
rect -581 -3459 -547 -3425
rect -917 -3527 -883 -3493
rect -849 -3527 -815 -3493
rect -649 -3527 -615 -3493
rect -581 -3527 -547 -3493
rect -97 -3191 -63 -3157
rect -29 -3191 5 -3157
rect 171 -3191 205 -3157
rect 239 -3191 273 -3157
rect -97 -3259 -63 -3225
rect 239 -3259 273 -3225
rect -97 -3459 -63 -3425
rect 239 -3459 273 -3425
rect -97 -3527 -63 -3493
rect -29 -3527 5 -3493
rect 171 -3527 205 -3493
rect 239 -3527 273 -3493
rect 723 -3191 757 -3157
rect 791 -3191 825 -3157
rect 991 -3191 1025 -3157
rect 1059 -3191 1093 -3157
rect 723 -3259 757 -3225
rect 1059 -3259 1093 -3225
rect 723 -3459 757 -3425
rect 1059 -3459 1093 -3425
rect 723 -3527 757 -3493
rect 791 -3527 825 -3493
rect 991 -3527 1025 -3493
rect 1059 -3527 1093 -3493
rect 1543 -3191 1577 -3157
rect 1611 -3191 1645 -3157
rect 1811 -3191 1845 -3157
rect 1879 -3191 1913 -3157
rect 1543 -3259 1577 -3225
rect 1879 -3259 1913 -3225
rect 1543 -3459 1577 -3425
rect 1879 -3459 1913 -3425
rect 1543 -3527 1577 -3493
rect 1611 -3527 1645 -3493
rect 1811 -3527 1845 -3493
rect 1879 -3527 1913 -3493
rect 2363 -3191 2397 -3157
rect 2431 -3191 2465 -3157
rect 2631 -3191 2665 -3157
rect 2699 -3191 2733 -3157
rect 2363 -3259 2397 -3225
rect 2699 -3259 2733 -3225
rect 2363 -3459 2397 -3425
rect 2699 -3459 2733 -3425
rect 2363 -3527 2397 -3493
rect 2431 -3527 2465 -3493
rect 2631 -3527 2665 -3493
rect 2699 -3527 2733 -3493
rect 3183 -3191 3217 -3157
rect 3251 -3191 3285 -3157
rect 3451 -3191 3485 -3157
rect 3519 -3191 3553 -3157
rect 3183 -3259 3217 -3225
rect 3519 -3259 3553 -3225
rect 3183 -3459 3217 -3425
rect 3519 -3459 3553 -3425
rect 3183 -3527 3217 -3493
rect 3251 -3527 3285 -3493
rect 3451 -3527 3485 -3493
rect 3519 -3527 3553 -3493
rect 4003 -3191 4037 -3157
rect 4071 -3191 4105 -3157
rect 4271 -3191 4305 -3157
rect 4339 -3191 4373 -3157
rect 4003 -3259 4037 -3225
rect 4339 -3259 4373 -3225
rect 4003 -3459 4037 -3425
rect 4339 -3459 4373 -3425
rect 4003 -3527 4037 -3493
rect 4071 -3527 4105 -3493
rect 4271 -3527 4305 -3493
rect 4339 -3527 4373 -3493
rect 4823 -3191 4857 -3157
rect 4891 -3191 4925 -3157
rect 5091 -3191 5125 -3157
rect 5159 -3191 5193 -3157
rect 4823 -3259 4857 -3225
rect 5159 -3259 5193 -3225
rect 4823 -3459 4857 -3425
rect 5159 -3459 5193 -3425
rect 4823 -3527 4857 -3493
rect 4891 -3527 4925 -3493
rect 5091 -3527 5125 -3493
rect 5159 -3527 5193 -3493
rect 5643 -3191 5677 -3157
rect 5711 -3191 5745 -3157
rect 5911 -3191 5945 -3157
rect 5979 -3191 6013 -3157
rect 5643 -3259 5677 -3225
rect 5979 -3259 6013 -3225
rect 5643 -3459 5677 -3425
rect 5979 -3459 6013 -3425
rect 5643 -3527 5677 -3493
rect 5711 -3527 5745 -3493
rect 5911 -3527 5945 -3493
rect 5979 -3527 6013 -3493
rect 6463 -3191 6497 -3157
rect 6531 -3191 6565 -3157
rect 6731 -3191 6765 -3157
rect 6799 -3191 6833 -3157
rect 6463 -3259 6497 -3225
rect 6799 -3259 6833 -3225
rect 6463 -3459 6497 -3425
rect 6799 -3459 6833 -3425
rect 6463 -3527 6497 -3493
rect 6531 -3527 6565 -3493
rect 6731 -3527 6765 -3493
rect 6799 -3527 6833 -3493
rect -917 -4011 -883 -3977
rect -849 -4011 -815 -3977
rect -649 -4011 -615 -3977
rect -581 -4011 -547 -3977
rect -917 -4079 -883 -4045
rect -581 -4079 -547 -4045
rect -917 -4279 -883 -4245
rect -581 -4279 -547 -4245
rect -917 -4347 -883 -4313
rect -849 -4347 -815 -4313
rect -649 -4347 -615 -4313
rect -581 -4347 -547 -4313
rect -97 -4011 -63 -3977
rect -29 -4011 5 -3977
rect 171 -4011 205 -3977
rect 239 -4011 273 -3977
rect -97 -4079 -63 -4045
rect 239 -4079 273 -4045
rect -97 -4279 -63 -4245
rect 239 -4279 273 -4245
rect -97 -4347 -63 -4313
rect -29 -4347 5 -4313
rect 171 -4347 205 -4313
rect 239 -4347 273 -4313
rect 723 -4011 757 -3977
rect 791 -4011 825 -3977
rect 991 -4011 1025 -3977
rect 1059 -4011 1093 -3977
rect 723 -4079 757 -4045
rect 1059 -4079 1093 -4045
rect 723 -4279 757 -4245
rect 1059 -4279 1093 -4245
rect 723 -4347 757 -4313
rect 791 -4347 825 -4313
rect 991 -4347 1025 -4313
rect 1059 -4347 1093 -4313
rect 1543 -4011 1577 -3977
rect 1611 -4011 1645 -3977
rect 1811 -4011 1845 -3977
rect 1879 -4011 1913 -3977
rect 1543 -4079 1577 -4045
rect 1879 -4079 1913 -4045
rect 1543 -4279 1577 -4245
rect 1879 -4279 1913 -4245
rect 1543 -4347 1577 -4313
rect 1611 -4347 1645 -4313
rect 1811 -4347 1845 -4313
rect 1879 -4347 1913 -4313
rect 2363 -4011 2397 -3977
rect 2431 -4011 2465 -3977
rect 2631 -4011 2665 -3977
rect 2699 -4011 2733 -3977
rect 2363 -4079 2397 -4045
rect 2699 -4079 2733 -4045
rect 2363 -4279 2397 -4245
rect 2699 -4279 2733 -4245
rect 2363 -4347 2397 -4313
rect 2431 -4347 2465 -4313
rect 2631 -4347 2665 -4313
rect 2699 -4347 2733 -4313
rect 3183 -4011 3217 -3977
rect 3251 -4011 3285 -3977
rect 3451 -4011 3485 -3977
rect 3519 -4011 3553 -3977
rect 3183 -4079 3217 -4045
rect 3519 -4079 3553 -4045
rect 3183 -4279 3217 -4245
rect 3519 -4279 3553 -4245
rect 3183 -4347 3217 -4313
rect 3251 -4347 3285 -4313
rect 3451 -4347 3485 -4313
rect 3519 -4347 3553 -4313
rect 4003 -4011 4037 -3977
rect 4071 -4011 4105 -3977
rect 4271 -4011 4305 -3977
rect 4339 -4011 4373 -3977
rect 4003 -4079 4037 -4045
rect 4339 -4079 4373 -4045
rect 4003 -4279 4037 -4245
rect 4339 -4279 4373 -4245
rect 4003 -4347 4037 -4313
rect 4071 -4347 4105 -4313
rect 4271 -4347 4305 -4313
rect 4339 -4347 4373 -4313
rect 4823 -4011 4857 -3977
rect 4891 -4011 4925 -3977
rect 5091 -4011 5125 -3977
rect 5159 -4011 5193 -3977
rect 4823 -4079 4857 -4045
rect 5159 -4079 5193 -4045
rect 4823 -4279 4857 -4245
rect 5159 -4279 5193 -4245
rect 4823 -4347 4857 -4313
rect 4891 -4347 4925 -4313
rect 5091 -4347 5125 -4313
rect 5159 -4347 5193 -4313
rect 5643 -4011 5677 -3977
rect 5711 -4011 5745 -3977
rect 5911 -4011 5945 -3977
rect 5979 -4011 6013 -3977
rect 5643 -4079 5677 -4045
rect 5979 -4079 6013 -4045
rect 5643 -4279 5677 -4245
rect 5979 -4279 6013 -4245
rect 5643 -4347 5677 -4313
rect 5711 -4347 5745 -4313
rect 5911 -4347 5945 -4313
rect 5979 -4347 6013 -4313
rect 6463 -4011 6497 -3977
rect 6531 -4011 6565 -3977
rect 6731 -4011 6765 -3977
rect 6799 -4011 6833 -3977
rect 6463 -4079 6497 -4045
rect 6799 -4079 6833 -4045
rect 6463 -4279 6497 -4245
rect 6799 -4279 6833 -4245
rect 6463 -4347 6497 -4313
rect 6531 -4347 6565 -4313
rect 6731 -4347 6765 -4313
rect 6799 -4347 6833 -4313
<< poly >>
rect 7500 6270 7530 6300
rect 7830 6270 7860 6300
rect 7500 4210 7530 4270
rect 7830 4210 7860 4270
rect 7480 4190 7560 4210
rect 7480 4150 7500 4190
rect 7540 4150 7560 4190
rect 7480 4130 7560 4150
rect 7800 4190 7880 4210
rect 7800 4150 7820 4190
rect 7860 4150 7880 4190
rect 7800 4130 7880 4150
rect 7500 4060 7530 4130
rect 7830 4060 7860 4130
rect 7500 2030 7530 2060
rect 7830 2030 7860 2060
<< polycont >>
rect 7500 4150 7540 4190
rect 7820 4150 7860 4190
<< xpolycontact >>
rect 8840 2800 9280 2940
rect 12080 2800 12520 2940
rect 15710 2800 16150 2940
rect 17000 2800 17440 2940
rect 6620 1300 6760 1740
rect 6620 10 6760 450
rect 7010 1300 7150 1740
rect 7010 10 7150 450
rect 7400 1300 7540 1740
rect 7400 10 7540 450
rect 7820 1300 7960 1740
rect 7820 10 7960 450
rect 15800 -1340 15940 -900
rect 15800 -3180 15940 -2740
rect 16190 -1340 16330 -900
rect 16190 -3180 16330 -2740
rect 16580 -1340 16720 -900
rect 16580 -3180 16720 -2740
rect 16970 -1340 17110 -900
rect 16970 -3180 17110 -2740
<< ppolyres >>
rect 9280 2800 12080 2940
rect 16150 2800 17000 2940
rect 6620 450 6760 1300
rect 7010 450 7150 1300
rect 7400 450 7540 1300
rect 7820 450 7960 1300
rect 15800 -2740 15940 -1340
rect 16190 -2740 16330 -1340
rect 16580 -2740 16720 -1340
rect 16970 -2740 17110 -1340
<< locali >>
rect 7400 6240 7490 6260
rect 6700 4400 6780 4420
rect 6700 4360 6720 4400
rect 6760 4360 6780 4400
rect 6700 1740 6780 4360
rect 7400 4300 7430 6240
rect 7470 4300 7490 6240
rect 7400 4250 7490 4300
rect 7540 6240 7820 6260
rect 7540 4300 7560 6240
rect 7600 4300 7660 6240
rect 7700 4300 7760 6240
rect 7800 4300 7820 6240
rect 7540 4250 7820 4300
rect 7870 6240 7960 6260
rect 7870 4300 7890 6240
rect 7930 4710 7960 6240
rect 7930 4690 8130 4710
rect 7930 4650 8070 4690
rect 8110 4650 8130 4690
rect 7930 4630 8130 4650
rect 7930 4300 7960 4630
rect 7870 4250 7960 4300
rect 7400 4090 7440 4250
rect 7480 4190 7560 4210
rect 7480 4150 7500 4190
rect 7540 4150 7560 4190
rect 7480 4130 7560 4150
rect 7600 4090 7760 4250
rect 7800 4190 7880 4210
rect 7800 4150 7820 4190
rect 7860 4150 7880 4190
rect 7800 4130 7880 4150
rect 7920 4090 7960 4250
rect 7400 4030 7490 4090
rect 7240 3960 7320 3980
rect 7240 3920 7260 3960
rect 7300 3920 7320 3960
rect 6760 1300 7010 1740
rect 7240 610 7320 3920
rect 7400 2090 7430 4030
rect 7470 2090 7490 4030
rect 7400 1740 7490 2090
rect 7540 4030 7820 4090
rect 7540 2090 7560 4030
rect 7600 2090 7660 4030
rect 7700 2090 7760 4030
rect 7800 2090 7820 4030
rect 7540 2070 7820 2090
rect 7870 4030 7960 4090
rect 7870 2090 7890 4030
rect 7930 2090 7960 4030
rect 8590 2910 8840 2940
rect 8590 2830 8650 2910
rect 8730 2830 8840 2910
rect 8590 2800 8840 2830
rect 7870 1740 7960 2090
rect 15860 1260 15940 2800
rect 15860 1220 15880 1260
rect 15920 1220 15940 1260
rect 15860 1200 15940 1220
rect 15830 930 15940 950
rect 15830 780 15850 930
rect 15920 780 15940 930
rect 7240 570 7260 610
rect 7300 570 7320 610
rect 7240 550 7320 570
rect 7650 610 7730 630
rect 7650 570 7670 610
rect 7710 570 7730 610
rect 7650 450 7730 570
rect 7150 10 7400 450
rect 7650 370 7820 450
rect 15830 260 15940 780
rect -1110 -544 7870 -510
rect -1110 -578 -1070 -544
rect -1036 -578 -1002 -544
rect -968 -578 -934 -544
rect -900 -578 -866 -544
rect -832 -578 -632 -544
rect -598 -578 -564 -544
rect -530 -578 -496 -544
rect -462 -578 -428 -544
rect -394 -578 -250 -544
rect -216 -578 -182 -544
rect -148 -578 -114 -544
rect -80 -578 -46 -544
rect -12 -578 188 -544
rect 222 -578 256 -544
rect 290 -578 324 -544
rect 358 -578 392 -544
rect 426 -578 570 -544
rect 604 -578 638 -544
rect 672 -578 706 -544
rect 740 -578 774 -544
rect 808 -578 1008 -544
rect 1042 -578 1076 -544
rect 1110 -578 1144 -544
rect 1178 -578 1212 -544
rect 1246 -578 1390 -544
rect 1424 -578 1458 -544
rect 1492 -578 1526 -544
rect 1560 -578 1594 -544
rect 1628 -578 1828 -544
rect 1862 -578 1896 -544
rect 1930 -578 1964 -544
rect 1998 -578 2032 -544
rect 2066 -578 2210 -544
rect 2244 -578 2278 -544
rect 2312 -578 2346 -544
rect 2380 -578 2414 -544
rect 2448 -578 2648 -544
rect 2682 -578 2716 -544
rect 2750 -578 2784 -544
rect 2818 -578 2852 -544
rect 2886 -578 3030 -544
rect 3064 -578 3098 -544
rect 3132 -578 3166 -544
rect 3200 -578 3234 -544
rect 3268 -578 3468 -544
rect 3502 -578 3536 -544
rect 3570 -578 3604 -544
rect 3638 -578 3672 -544
rect 3706 -578 3850 -544
rect 3884 -578 3918 -544
rect 3952 -578 3986 -544
rect 4020 -578 4054 -544
rect 4088 -578 4288 -544
rect 4322 -578 4356 -544
rect 4390 -578 4424 -544
rect 4458 -578 4492 -544
rect 4526 -578 4670 -544
rect 4704 -578 4738 -544
rect 4772 -578 4806 -544
rect 4840 -578 4874 -544
rect 4908 -578 5108 -544
rect 5142 -578 5176 -544
rect 5210 -578 5244 -544
rect 5278 -578 5312 -544
rect 5346 -578 5490 -544
rect 5524 -578 5558 -544
rect 5592 -578 5626 -544
rect 5660 -578 5694 -544
rect 5728 -578 5928 -544
rect 5962 -578 5996 -544
rect 6030 -578 6064 -544
rect 6098 -578 6132 -544
rect 6166 -578 6310 -544
rect 6344 -578 6378 -544
rect 6412 -578 6446 -544
rect 6480 -578 6514 -544
rect 6548 -578 6748 -544
rect 6782 -578 6816 -544
rect 6850 -578 6884 -544
rect 6918 -578 6952 -544
rect 6986 -578 7160 -544
rect 7194 -578 7228 -544
rect 7262 -578 7296 -544
rect 7330 -578 7364 -544
rect 7398 -578 7598 -544
rect 7632 -578 7666 -544
rect 7700 -578 7734 -544
rect 7768 -578 7802 -544
rect 7836 -578 7870 -544
rect -1110 -611 7870 -578
rect -1110 -612 7360 -611
rect -1110 -646 -1070 -612
rect -1036 -646 -428 -612
rect -394 -646 -250 -612
rect -216 -646 392 -612
rect 426 -646 570 -612
rect 604 -646 1212 -612
rect 1246 -646 1390 -612
rect 1424 -646 2032 -612
rect 2066 -646 2210 -612
rect 2244 -646 2852 -612
rect 2886 -646 3030 -612
rect 3064 -646 3672 -612
rect 3706 -646 3850 -612
rect 3884 -646 4492 -612
rect 4526 -646 4670 -612
rect 4704 -646 5312 -612
rect 5346 -646 5490 -612
rect 5524 -646 6132 -612
rect 6166 -646 6310 -612
rect 6344 -646 6952 -612
rect 6986 -646 7160 -612
rect 7194 -646 7360 -612
rect -1110 -673 7360 -646
rect 7769 -612 7870 -611
rect 7769 -646 7802 -612
rect 7836 -646 7870 -612
rect -1110 -680 7707 -673
rect -1110 -714 -1070 -680
rect -1036 -697 -428 -680
rect -1036 -714 -917 -697
rect -1110 -731 -917 -714
rect -883 -731 -849 -697
rect -815 -731 -649 -697
rect -615 -731 -581 -697
rect -547 -714 -428 -697
rect -394 -714 -250 -680
rect -216 -697 392 -680
rect -216 -714 -97 -697
rect -547 -731 -97 -714
rect -63 -731 -29 -697
rect 5 -731 171 -697
rect 205 -731 239 -697
rect 273 -714 392 -697
rect 426 -714 570 -680
rect 604 -697 1212 -680
rect 604 -714 723 -697
rect 273 -731 723 -714
rect 757 -731 791 -697
rect 825 -731 991 -697
rect 1025 -731 1059 -697
rect 1093 -714 1212 -697
rect 1246 -714 1390 -680
rect 1424 -697 2032 -680
rect 1424 -714 1543 -697
rect 1093 -731 1543 -714
rect 1577 -731 1611 -697
rect 1645 -731 1811 -697
rect 1845 -731 1879 -697
rect 1913 -714 2032 -697
rect 2066 -714 2210 -680
rect 2244 -697 2852 -680
rect 2244 -714 2363 -697
rect 1913 -731 2363 -714
rect 2397 -731 2431 -697
rect 2465 -731 2631 -697
rect 2665 -731 2699 -697
rect 2733 -714 2852 -697
rect 2886 -714 3030 -680
rect 3064 -697 3672 -680
rect 3064 -714 3183 -697
rect 2733 -731 3183 -714
rect 3217 -731 3251 -697
rect 3285 -731 3451 -697
rect 3485 -731 3519 -697
rect 3553 -714 3672 -697
rect 3706 -714 3850 -680
rect 3884 -697 4492 -680
rect 3884 -714 4003 -697
rect 3553 -731 4003 -714
rect 4037 -731 4071 -697
rect 4105 -731 4271 -697
rect 4305 -731 4339 -697
rect 4373 -714 4492 -697
rect 4526 -714 4670 -680
rect 4704 -697 5312 -680
rect 4704 -714 4823 -697
rect 4373 -731 4823 -714
rect 4857 -731 4891 -697
rect 4925 -731 5091 -697
rect 5125 -731 5159 -697
rect 5193 -714 5312 -697
rect 5346 -714 5490 -680
rect 5524 -697 6132 -680
rect 5524 -714 5643 -697
rect 5193 -731 5643 -714
rect 5677 -731 5711 -697
rect 5745 -731 5911 -697
rect 5945 -731 5979 -697
rect 6013 -714 6132 -697
rect 6166 -714 6310 -680
rect 6344 -697 6952 -680
rect 6344 -714 6463 -697
rect 6013 -731 6463 -714
rect 6497 -731 6531 -697
rect 6565 -731 6731 -697
rect 6765 -731 6799 -697
rect 6833 -714 6952 -697
rect 6986 -714 7160 -680
rect 7194 -697 7707 -680
rect 7194 -714 7313 -697
rect 6833 -731 7313 -714
rect 7347 -731 7381 -697
rect 7415 -731 7581 -697
rect 7615 -731 7649 -697
rect 7683 -731 7707 -697
rect -1110 -745 7707 -731
rect -1110 -748 7361 -745
rect -1110 -750 -1070 -748
rect -1104 -782 -1070 -750
rect -1036 -750 -428 -748
rect -1036 -782 -1003 -750
rect -1104 -982 -1003 -782
rect -1104 -1010 -1070 -982
rect -1110 -1016 -1070 -1010
rect -1036 -1010 -1003 -982
rect -941 -765 -869 -750
rect -941 -799 -917 -765
rect -883 -799 -869 -765
rect -941 -965 -869 -799
rect -595 -765 -523 -750
rect -595 -799 -581 -765
rect -547 -799 -523 -765
rect -811 -817 -653 -803
rect -811 -851 -797 -817
rect -763 -831 -701 -817
rect -667 -851 -653 -817
rect -811 -913 -783 -851
rect -681 -913 -653 -851
rect -811 -947 -797 -913
rect -763 -947 -701 -933
rect -667 -947 -653 -913
rect -811 -961 -653 -947
rect -941 -999 -917 -965
rect -883 -999 -869 -965
rect -941 -1010 -869 -999
rect -595 -965 -523 -799
rect -595 -999 -581 -965
rect -547 -999 -523 -965
rect -595 -1010 -523 -999
rect -461 -782 -428 -750
rect -394 -750 -250 -748
rect -394 -782 -360 -750
rect -461 -982 -360 -782
rect -461 -1010 -428 -982
rect -1036 -1016 -428 -1010
rect -394 -1010 -360 -982
rect -284 -782 -250 -750
rect -216 -750 392 -748
rect -216 -782 -183 -750
rect -284 -982 -183 -782
rect -284 -1010 -250 -982
rect -394 -1016 -250 -1010
rect -216 -1010 -183 -982
rect -121 -765 -49 -750
rect -121 -799 -97 -765
rect -63 -799 -49 -765
rect -121 -965 -49 -799
rect 225 -765 297 -750
rect 225 -799 239 -765
rect 273 -799 297 -765
rect 9 -817 167 -803
rect 9 -851 23 -817
rect 57 -831 119 -817
rect 153 -851 167 -817
rect 9 -913 37 -851
rect 139 -913 167 -851
rect 9 -947 23 -913
rect 57 -947 119 -933
rect 153 -947 167 -913
rect 9 -961 167 -947
rect -121 -999 -97 -965
rect -63 -999 -49 -965
rect -121 -1010 -49 -999
rect 225 -965 297 -799
rect 225 -999 239 -965
rect 273 -999 297 -965
rect 225 -1010 297 -999
rect 359 -782 392 -750
rect 426 -750 570 -748
rect 426 -782 460 -750
rect 359 -982 460 -782
rect 359 -1010 392 -982
rect -216 -1016 392 -1010
rect 426 -1010 460 -982
rect 536 -782 570 -750
rect 604 -750 1212 -748
rect 604 -782 637 -750
rect 536 -982 637 -782
rect 536 -1010 570 -982
rect 426 -1016 570 -1010
rect 604 -1010 637 -982
rect 699 -765 771 -750
rect 699 -799 723 -765
rect 757 -799 771 -765
rect 699 -965 771 -799
rect 1045 -765 1117 -750
rect 1045 -799 1059 -765
rect 1093 -799 1117 -765
rect 829 -817 987 -803
rect 829 -851 843 -817
rect 877 -831 939 -817
rect 973 -851 987 -817
rect 829 -913 857 -851
rect 959 -913 987 -851
rect 829 -947 843 -913
rect 877 -947 939 -933
rect 973 -947 987 -913
rect 829 -961 987 -947
rect 699 -999 723 -965
rect 757 -999 771 -965
rect 699 -1010 771 -999
rect 1045 -965 1117 -799
rect 1045 -999 1059 -965
rect 1093 -999 1117 -965
rect 1045 -1010 1117 -999
rect 1179 -782 1212 -750
rect 1246 -750 1390 -748
rect 1246 -782 1280 -750
rect 1179 -982 1280 -782
rect 1179 -1010 1212 -982
rect 604 -1016 1212 -1010
rect 1246 -1010 1280 -982
rect 1356 -782 1390 -750
rect 1424 -750 2032 -748
rect 1424 -782 1457 -750
rect 1356 -982 1457 -782
rect 1356 -1010 1390 -982
rect 1246 -1016 1390 -1010
rect 1424 -1010 1457 -982
rect 1519 -765 1591 -750
rect 1519 -799 1543 -765
rect 1577 -799 1591 -765
rect 1519 -965 1591 -799
rect 1865 -765 1937 -750
rect 1865 -799 1879 -765
rect 1913 -799 1937 -765
rect 1649 -817 1807 -803
rect 1649 -851 1663 -817
rect 1697 -831 1759 -817
rect 1793 -851 1807 -817
rect 1649 -913 1677 -851
rect 1779 -913 1807 -851
rect 1649 -947 1663 -913
rect 1697 -947 1759 -933
rect 1793 -947 1807 -913
rect 1649 -961 1807 -947
rect 1519 -999 1543 -965
rect 1577 -999 1591 -965
rect 1519 -1010 1591 -999
rect 1865 -965 1937 -799
rect 1865 -999 1879 -965
rect 1913 -999 1937 -965
rect 1865 -1010 1937 -999
rect 1999 -782 2032 -750
rect 2066 -750 2210 -748
rect 2066 -782 2100 -750
rect 1999 -982 2100 -782
rect 1999 -1010 2032 -982
rect 1424 -1016 2032 -1010
rect 2066 -1010 2100 -982
rect 2176 -782 2210 -750
rect 2244 -750 2852 -748
rect 2244 -782 2277 -750
rect 2176 -982 2277 -782
rect 2176 -1010 2210 -982
rect 2066 -1016 2210 -1010
rect 2244 -1010 2277 -982
rect 2339 -765 2411 -750
rect 2339 -799 2363 -765
rect 2397 -799 2411 -765
rect 2339 -965 2411 -799
rect 2685 -765 2757 -750
rect 2685 -799 2699 -765
rect 2733 -799 2757 -765
rect 2469 -817 2627 -803
rect 2469 -851 2483 -817
rect 2517 -831 2579 -817
rect 2613 -851 2627 -817
rect 2469 -913 2497 -851
rect 2599 -913 2627 -851
rect 2469 -947 2483 -913
rect 2517 -947 2579 -933
rect 2613 -947 2627 -913
rect 2469 -961 2627 -947
rect 2339 -999 2363 -965
rect 2397 -999 2411 -965
rect 2339 -1010 2411 -999
rect 2685 -965 2757 -799
rect 2685 -999 2699 -965
rect 2733 -999 2757 -965
rect 2685 -1010 2757 -999
rect 2819 -782 2852 -750
rect 2886 -750 3030 -748
rect 2886 -782 2920 -750
rect 2819 -982 2920 -782
rect 2819 -1010 2852 -982
rect 2244 -1016 2852 -1010
rect 2886 -1010 2920 -982
rect 2996 -782 3030 -750
rect 3064 -750 3672 -748
rect 3064 -782 3097 -750
rect 2996 -982 3097 -782
rect 2996 -1010 3030 -982
rect 2886 -1016 3030 -1010
rect 3064 -1010 3097 -982
rect 3159 -765 3231 -750
rect 3159 -799 3183 -765
rect 3217 -799 3231 -765
rect 3159 -965 3231 -799
rect 3505 -765 3577 -750
rect 3505 -799 3519 -765
rect 3553 -799 3577 -765
rect 3289 -817 3447 -803
rect 3289 -851 3303 -817
rect 3337 -831 3399 -817
rect 3433 -851 3447 -817
rect 3289 -913 3317 -851
rect 3419 -913 3447 -851
rect 3289 -947 3303 -913
rect 3337 -947 3399 -933
rect 3433 -947 3447 -913
rect 3289 -961 3447 -947
rect 3159 -999 3183 -965
rect 3217 -999 3231 -965
rect 3159 -1010 3231 -999
rect 3505 -965 3577 -799
rect 3505 -999 3519 -965
rect 3553 -999 3577 -965
rect 3505 -1010 3577 -999
rect 3639 -782 3672 -750
rect 3706 -750 3850 -748
rect 3706 -782 3740 -750
rect 3639 -982 3740 -782
rect 3639 -1010 3672 -982
rect 3064 -1016 3672 -1010
rect 3706 -1010 3740 -982
rect 3816 -782 3850 -750
rect 3884 -750 4492 -748
rect 3884 -782 3917 -750
rect 3816 -982 3917 -782
rect 3816 -1010 3850 -982
rect 3706 -1016 3850 -1010
rect 3884 -1010 3917 -982
rect 3979 -765 4051 -750
rect 3979 -799 4003 -765
rect 4037 -799 4051 -765
rect 3979 -965 4051 -799
rect 4325 -765 4397 -750
rect 4325 -799 4339 -765
rect 4373 -799 4397 -765
rect 4109 -817 4267 -803
rect 4109 -851 4123 -817
rect 4157 -831 4219 -817
rect 4253 -851 4267 -817
rect 4109 -913 4137 -851
rect 4239 -913 4267 -851
rect 4109 -947 4123 -913
rect 4157 -947 4219 -933
rect 4253 -947 4267 -913
rect 4109 -961 4267 -947
rect 3979 -999 4003 -965
rect 4037 -999 4051 -965
rect 3979 -1010 4051 -999
rect 4325 -965 4397 -799
rect 4325 -999 4339 -965
rect 4373 -999 4397 -965
rect 4325 -1010 4397 -999
rect 4459 -782 4492 -750
rect 4526 -750 4670 -748
rect 4526 -782 4560 -750
rect 4459 -982 4560 -782
rect 4459 -1010 4492 -982
rect 3884 -1016 4492 -1010
rect 4526 -1010 4560 -982
rect 4636 -782 4670 -750
rect 4704 -750 5312 -748
rect 4704 -782 4737 -750
rect 4636 -982 4737 -782
rect 4636 -1010 4670 -982
rect 4526 -1016 4670 -1010
rect 4704 -1010 4737 -982
rect 4799 -765 4871 -750
rect 4799 -799 4823 -765
rect 4857 -799 4871 -765
rect 4799 -965 4871 -799
rect 5145 -765 5217 -750
rect 5145 -799 5159 -765
rect 5193 -799 5217 -765
rect 4929 -817 5087 -803
rect 4929 -851 4943 -817
rect 4977 -831 5039 -817
rect 5073 -851 5087 -817
rect 4929 -913 4957 -851
rect 5059 -913 5087 -851
rect 4929 -947 4943 -913
rect 4977 -947 5039 -933
rect 5073 -947 5087 -913
rect 4929 -961 5087 -947
rect 4799 -999 4823 -965
rect 4857 -999 4871 -965
rect 4799 -1010 4871 -999
rect 5145 -965 5217 -799
rect 5145 -999 5159 -965
rect 5193 -999 5217 -965
rect 5145 -1010 5217 -999
rect 5279 -782 5312 -750
rect 5346 -750 5490 -748
rect 5346 -782 5380 -750
rect 5279 -982 5380 -782
rect 5279 -1010 5312 -982
rect 4704 -1016 5312 -1010
rect 5346 -1010 5380 -982
rect 5456 -782 5490 -750
rect 5524 -750 6132 -748
rect 5524 -782 5557 -750
rect 5456 -982 5557 -782
rect 5456 -1010 5490 -982
rect 5346 -1016 5490 -1010
rect 5524 -1010 5557 -982
rect 5619 -765 5691 -750
rect 5619 -799 5643 -765
rect 5677 -799 5691 -765
rect 5619 -965 5691 -799
rect 5965 -765 6037 -750
rect 5965 -799 5979 -765
rect 6013 -799 6037 -765
rect 5749 -817 5907 -803
rect 5749 -851 5763 -817
rect 5797 -831 5859 -817
rect 5893 -851 5907 -817
rect 5749 -913 5777 -851
rect 5879 -913 5907 -851
rect 5749 -947 5763 -913
rect 5797 -947 5859 -933
rect 5893 -947 5907 -913
rect 5749 -961 5907 -947
rect 5619 -999 5643 -965
rect 5677 -999 5691 -965
rect 5619 -1010 5691 -999
rect 5965 -965 6037 -799
rect 5965 -999 5979 -965
rect 6013 -999 6037 -965
rect 5965 -1010 6037 -999
rect 6099 -782 6132 -750
rect 6166 -750 6310 -748
rect 6166 -782 6200 -750
rect 6099 -982 6200 -782
rect 6099 -1010 6132 -982
rect 5524 -1016 6132 -1010
rect 6166 -1010 6200 -982
rect 6276 -782 6310 -750
rect 6344 -750 6952 -748
rect 6344 -782 6377 -750
rect 6276 -982 6377 -782
rect 6276 -1010 6310 -982
rect 6166 -1016 6310 -1010
rect 6344 -1010 6377 -982
rect 6439 -765 6511 -750
rect 6439 -799 6463 -765
rect 6497 -799 6511 -765
rect 6439 -965 6511 -799
rect 6785 -765 6857 -750
rect 6785 -799 6799 -765
rect 6833 -799 6857 -765
rect 6569 -817 6727 -803
rect 6569 -851 6583 -817
rect 6617 -831 6679 -817
rect 6713 -851 6727 -817
rect 6569 -913 6597 -851
rect 6699 -913 6727 -851
rect 6569 -947 6583 -913
rect 6617 -947 6679 -933
rect 6713 -947 6727 -913
rect 6569 -961 6727 -947
rect 6439 -999 6463 -965
rect 6497 -999 6511 -965
rect 6439 -1010 6511 -999
rect 6785 -965 6857 -799
rect 6785 -999 6799 -965
rect 6833 -999 6857 -965
rect 6785 -1010 6857 -999
rect 6919 -782 6952 -750
rect 6986 -782 7160 -748
rect 7194 -765 7361 -748
rect 7194 -782 7313 -765
rect 6919 -799 7313 -782
rect 7347 -799 7361 -765
rect 6919 -965 7361 -799
rect 7635 -765 7707 -745
rect 7635 -799 7649 -765
rect 7683 -799 7707 -765
rect 7419 -817 7577 -803
rect 7419 -851 7433 -817
rect 7467 -831 7529 -817
rect 7563 -851 7577 -817
rect 7419 -913 7447 -851
rect 7549 -913 7577 -851
rect 7419 -947 7433 -913
rect 7467 -947 7529 -933
rect 7563 -947 7577 -913
rect 7419 -961 7577 -947
rect 6919 -982 7313 -965
rect 6919 -1010 6952 -982
rect 6344 -1016 6952 -1010
rect 6986 -1016 7160 -982
rect 7194 -999 7313 -982
rect 7347 -999 7361 -965
rect 7194 -1016 7361 -999
rect -1110 -1019 7361 -1016
rect 7635 -965 7707 -799
rect 7635 -999 7649 -965
rect 7683 -999 7707 -965
rect 7635 -1019 7707 -999
rect -1110 -1033 7707 -1019
rect -1110 -1050 -917 -1033
rect -1110 -1084 -1070 -1050
rect -1036 -1067 -917 -1050
rect -883 -1067 -849 -1033
rect -815 -1067 -649 -1033
rect -615 -1067 -581 -1033
rect -547 -1050 -97 -1033
rect -547 -1067 -428 -1050
rect -1036 -1084 -428 -1067
rect -394 -1084 -250 -1050
rect -216 -1067 -97 -1050
rect -63 -1067 -29 -1033
rect 5 -1067 171 -1033
rect 205 -1067 239 -1033
rect 273 -1050 723 -1033
rect 273 -1067 392 -1050
rect -216 -1084 392 -1067
rect 426 -1084 570 -1050
rect 604 -1067 723 -1050
rect 757 -1067 791 -1033
rect 825 -1067 991 -1033
rect 1025 -1067 1059 -1033
rect 1093 -1050 1543 -1033
rect 1093 -1067 1212 -1050
rect 604 -1084 1212 -1067
rect 1246 -1084 1390 -1050
rect 1424 -1067 1543 -1050
rect 1577 -1067 1611 -1033
rect 1645 -1067 1811 -1033
rect 1845 -1067 1879 -1033
rect 1913 -1050 2363 -1033
rect 1913 -1067 2032 -1050
rect 1424 -1084 2032 -1067
rect 2066 -1084 2210 -1050
rect 2244 -1067 2363 -1050
rect 2397 -1067 2431 -1033
rect 2465 -1067 2631 -1033
rect 2665 -1067 2699 -1033
rect 2733 -1050 3183 -1033
rect 2733 -1067 2852 -1050
rect 2244 -1084 2852 -1067
rect 2886 -1084 3030 -1050
rect 3064 -1067 3183 -1050
rect 3217 -1067 3251 -1033
rect 3285 -1067 3451 -1033
rect 3485 -1067 3519 -1033
rect 3553 -1050 4003 -1033
rect 3553 -1067 3672 -1050
rect 3064 -1084 3672 -1067
rect 3706 -1084 3850 -1050
rect 3884 -1067 4003 -1050
rect 4037 -1067 4071 -1033
rect 4105 -1067 4271 -1033
rect 4305 -1067 4339 -1033
rect 4373 -1050 4823 -1033
rect 4373 -1067 4492 -1050
rect 3884 -1084 4492 -1067
rect 4526 -1084 4670 -1050
rect 4704 -1067 4823 -1050
rect 4857 -1067 4891 -1033
rect 4925 -1067 5091 -1033
rect 5125 -1067 5159 -1033
rect 5193 -1050 5643 -1033
rect 5193 -1067 5312 -1050
rect 4704 -1084 5312 -1067
rect 5346 -1084 5490 -1050
rect 5524 -1067 5643 -1050
rect 5677 -1067 5711 -1033
rect 5745 -1067 5911 -1033
rect 5945 -1067 5979 -1033
rect 6013 -1050 6463 -1033
rect 6013 -1067 6132 -1050
rect 5524 -1084 6132 -1067
rect 6166 -1084 6310 -1050
rect 6344 -1067 6463 -1050
rect 6497 -1067 6531 -1033
rect 6565 -1067 6731 -1033
rect 6765 -1067 6799 -1033
rect 6833 -1050 7313 -1033
rect 6833 -1067 6952 -1050
rect 6344 -1084 6952 -1067
rect 6986 -1084 7160 -1050
rect 7194 -1067 7313 -1050
rect 7347 -1067 7381 -1033
rect 7415 -1067 7581 -1033
rect 7615 -1067 7649 -1033
rect 7683 -1067 7707 -1033
rect 7194 -1084 7707 -1067
rect -1110 -1091 7707 -1084
rect 7769 -680 7870 -646
rect 7769 -714 7802 -680
rect 7836 -714 7870 -680
rect 7769 -748 7870 -714
rect 7769 -782 7802 -748
rect 7836 -782 7870 -748
rect 7769 -982 7870 -782
rect 7769 -1016 7802 -982
rect 7836 -1016 7870 -982
rect 7769 -1050 7870 -1016
rect 7769 -1084 7802 -1050
rect 7836 -1084 7870 -1050
rect -1110 -1118 7360 -1091
rect -1110 -1152 -1070 -1118
rect -1036 -1152 -428 -1118
rect -394 -1152 -250 -1118
rect -216 -1152 392 -1118
rect 426 -1152 570 -1118
rect 604 -1152 1212 -1118
rect 1246 -1152 1390 -1118
rect 1424 -1152 2032 -1118
rect 2066 -1152 2210 -1118
rect 2244 -1152 2852 -1118
rect 2886 -1152 3030 -1118
rect 3064 -1152 3672 -1118
rect 3706 -1152 3850 -1118
rect 3884 -1152 4492 -1118
rect 4526 -1152 4670 -1118
rect 4704 -1152 5312 -1118
rect 5346 -1152 5490 -1118
rect 5524 -1152 6132 -1118
rect 6166 -1152 6310 -1118
rect 6344 -1152 6952 -1118
rect 6986 -1152 7160 -1118
rect 7194 -1140 7360 -1118
rect 7769 -1118 7870 -1084
rect 7769 -1140 7802 -1118
rect 7194 -1152 7802 -1140
rect 7836 -1140 7870 -1118
rect 15800 -900 15940 260
rect 7836 -1152 8790 -1140
rect -1110 -1170 8790 -1152
rect -1110 -1186 8620 -1170
rect -1110 -1220 -1070 -1186
rect -1036 -1220 -1002 -1186
rect -968 -1220 -934 -1186
rect -900 -1220 -866 -1186
rect -832 -1220 -632 -1186
rect -598 -1220 -564 -1186
rect -530 -1220 -496 -1186
rect -462 -1220 -428 -1186
rect -394 -1220 -250 -1186
rect -216 -1220 -182 -1186
rect -148 -1220 -114 -1186
rect -80 -1220 -46 -1186
rect -12 -1220 188 -1186
rect 222 -1220 256 -1186
rect 290 -1220 324 -1186
rect 358 -1220 392 -1186
rect 426 -1220 570 -1186
rect 604 -1220 638 -1186
rect 672 -1220 706 -1186
rect 740 -1220 774 -1186
rect 808 -1220 1008 -1186
rect 1042 -1220 1076 -1186
rect 1110 -1220 1144 -1186
rect 1178 -1220 1212 -1186
rect 1246 -1220 1390 -1186
rect 1424 -1220 1458 -1186
rect 1492 -1220 1526 -1186
rect 1560 -1220 1594 -1186
rect 1628 -1220 1828 -1186
rect 1862 -1220 1896 -1186
rect 1930 -1220 1964 -1186
rect 1998 -1220 2032 -1186
rect 2066 -1220 2210 -1186
rect 2244 -1220 2278 -1186
rect 2312 -1220 2346 -1186
rect 2380 -1220 2414 -1186
rect 2448 -1220 2648 -1186
rect 2682 -1220 2716 -1186
rect 2750 -1220 2784 -1186
rect 2818 -1220 2852 -1186
rect 2886 -1220 3030 -1186
rect 3064 -1220 3098 -1186
rect 3132 -1220 3166 -1186
rect 3200 -1220 3234 -1186
rect 3268 -1220 3468 -1186
rect 3502 -1220 3536 -1186
rect 3570 -1220 3604 -1186
rect 3638 -1220 3672 -1186
rect 3706 -1220 3850 -1186
rect 3884 -1220 3918 -1186
rect 3952 -1220 3986 -1186
rect 4020 -1220 4054 -1186
rect 4088 -1220 4288 -1186
rect 4322 -1220 4356 -1186
rect 4390 -1220 4424 -1186
rect 4458 -1220 4492 -1186
rect 4526 -1220 4670 -1186
rect 4704 -1220 4738 -1186
rect 4772 -1220 4806 -1186
rect 4840 -1220 4874 -1186
rect 4908 -1220 5108 -1186
rect 5142 -1220 5176 -1186
rect 5210 -1220 5244 -1186
rect 5278 -1220 5312 -1186
rect 5346 -1220 5490 -1186
rect 5524 -1220 5558 -1186
rect 5592 -1220 5626 -1186
rect 5660 -1220 5694 -1186
rect 5728 -1220 5928 -1186
rect 5962 -1220 5996 -1186
rect 6030 -1220 6064 -1186
rect 6098 -1220 6132 -1186
rect 6166 -1220 6310 -1186
rect 6344 -1220 6378 -1186
rect 6412 -1220 6446 -1186
rect 6480 -1220 6514 -1186
rect 6548 -1220 6748 -1186
rect 6782 -1220 6816 -1186
rect 6850 -1220 6884 -1186
rect 6918 -1220 6952 -1186
rect 6986 -1220 7160 -1186
rect 7194 -1220 7228 -1186
rect 7262 -1220 7296 -1186
rect 7330 -1220 7364 -1186
rect 7398 -1220 7598 -1186
rect 7632 -1220 7666 -1186
rect 7700 -1220 7734 -1186
rect 7768 -1220 7802 -1186
rect 7836 -1220 8620 -1186
rect -1110 -1364 8620 -1220
rect -1110 -1398 -1070 -1364
rect -1036 -1398 -1002 -1364
rect -968 -1398 -934 -1364
rect -900 -1398 -866 -1364
rect -832 -1398 -632 -1364
rect -598 -1398 -564 -1364
rect -530 -1398 -496 -1364
rect -462 -1398 -428 -1364
rect -394 -1398 -250 -1364
rect -216 -1398 -182 -1364
rect -148 -1398 -114 -1364
rect -80 -1398 -46 -1364
rect -12 -1398 188 -1364
rect 222 -1398 256 -1364
rect 290 -1398 324 -1364
rect 358 -1398 392 -1364
rect 426 -1398 570 -1364
rect 604 -1398 638 -1364
rect 672 -1398 706 -1364
rect 740 -1398 774 -1364
rect 808 -1398 1008 -1364
rect 1042 -1398 1076 -1364
rect 1110 -1398 1144 -1364
rect 1178 -1398 1212 -1364
rect 1246 -1398 1390 -1364
rect 1424 -1398 1458 -1364
rect 1492 -1398 1526 -1364
rect 1560 -1398 1594 -1364
rect 1628 -1398 1828 -1364
rect 1862 -1398 1896 -1364
rect 1930 -1398 1964 -1364
rect 1998 -1398 2032 -1364
rect 2066 -1398 2210 -1364
rect 2244 -1398 2278 -1364
rect 2312 -1398 2346 -1364
rect 2380 -1398 2414 -1364
rect 2448 -1398 2648 -1364
rect 2682 -1398 2716 -1364
rect 2750 -1398 2784 -1364
rect 2818 -1398 2852 -1364
rect 2886 -1398 3030 -1364
rect 3064 -1398 3098 -1364
rect 3132 -1398 3166 -1364
rect 3200 -1398 3234 -1364
rect 3268 -1398 3468 -1364
rect 3502 -1398 3536 -1364
rect 3570 -1398 3604 -1364
rect 3638 -1398 3672 -1364
rect 3706 -1398 3850 -1364
rect 3884 -1398 3918 -1364
rect 3952 -1398 3986 -1364
rect 4020 -1398 4054 -1364
rect 4088 -1398 4288 -1364
rect 4322 -1398 4356 -1364
rect 4390 -1398 4424 -1364
rect 4458 -1398 4492 -1364
rect 4526 -1398 4670 -1364
rect 4704 -1398 4738 -1364
rect 4772 -1398 4806 -1364
rect 4840 -1398 4874 -1364
rect 4908 -1398 5108 -1364
rect 5142 -1398 5176 -1364
rect 5210 -1398 5244 -1364
rect 5278 -1398 5312 -1364
rect 5346 -1398 5490 -1364
rect 5524 -1398 5558 -1364
rect 5592 -1398 5626 -1364
rect 5660 -1398 5694 -1364
rect 5728 -1398 5928 -1364
rect 5962 -1398 5996 -1364
rect 6030 -1398 6064 -1364
rect 6098 -1398 6132 -1364
rect 6166 -1398 6310 -1364
rect 6344 -1398 6378 -1364
rect 6412 -1398 6446 -1364
rect 6480 -1398 6514 -1364
rect 6548 -1398 6748 -1364
rect 6782 -1398 6816 -1364
rect 6850 -1398 6884 -1364
rect 6918 -1398 6952 -1364
rect 6986 -1398 8620 -1364
rect -1110 -1432 8620 -1398
rect -1110 -1466 -1070 -1432
rect -1036 -1466 -428 -1432
rect -394 -1466 -250 -1432
rect -216 -1466 392 -1432
rect 426 -1466 570 -1432
rect 604 -1466 1212 -1432
rect 1246 -1466 1390 -1432
rect 1424 -1466 2032 -1432
rect 2066 -1466 2210 -1432
rect 2244 -1466 2852 -1432
rect 2886 -1466 3030 -1432
rect 3064 -1466 3672 -1432
rect 3706 -1466 3850 -1432
rect 3884 -1466 4492 -1432
rect 4526 -1466 4670 -1432
rect 4704 -1466 5312 -1432
rect 5346 -1466 5490 -1432
rect 5524 -1466 6132 -1432
rect 6166 -1466 6310 -1432
rect 6344 -1466 6952 -1432
rect 6986 -1466 8620 -1432
rect -1110 -1500 8620 -1466
rect -1110 -1534 -1070 -1500
rect -1036 -1517 -428 -1500
rect -1036 -1534 -917 -1517
rect -1110 -1551 -917 -1534
rect -883 -1551 -849 -1517
rect -815 -1551 -649 -1517
rect -615 -1551 -581 -1517
rect -547 -1534 -428 -1517
rect -394 -1534 -250 -1500
rect -216 -1517 392 -1500
rect -216 -1534 -97 -1517
rect -547 -1551 -97 -1534
rect -63 -1551 -29 -1517
rect 5 -1551 171 -1517
rect 205 -1551 239 -1517
rect 273 -1534 392 -1517
rect 426 -1534 570 -1500
rect 604 -1517 1212 -1500
rect 604 -1534 723 -1517
rect 273 -1551 723 -1534
rect 757 -1551 791 -1517
rect 825 -1551 991 -1517
rect 1025 -1551 1059 -1517
rect 1093 -1534 1212 -1517
rect 1246 -1534 1390 -1500
rect 1424 -1517 2032 -1500
rect 1424 -1534 1543 -1517
rect 1093 -1551 1543 -1534
rect 1577 -1551 1611 -1517
rect 1645 -1551 1811 -1517
rect 1845 -1551 1879 -1517
rect 1913 -1534 2032 -1517
rect 2066 -1534 2210 -1500
rect 2244 -1517 2852 -1500
rect 2244 -1534 2363 -1517
rect 1913 -1551 2363 -1534
rect 2397 -1551 2431 -1517
rect 2465 -1551 2631 -1517
rect 2665 -1551 2699 -1517
rect 2733 -1534 2852 -1517
rect 2886 -1534 3030 -1500
rect 3064 -1517 3672 -1500
rect 3064 -1534 3183 -1517
rect 2733 -1551 3183 -1534
rect 3217 -1551 3251 -1517
rect 3285 -1551 3451 -1517
rect 3485 -1551 3519 -1517
rect 3553 -1534 3672 -1517
rect 3706 -1534 3850 -1500
rect 3884 -1517 4492 -1500
rect 3884 -1534 4003 -1517
rect 3553 -1551 4003 -1534
rect 4037 -1551 4071 -1517
rect 4105 -1551 4271 -1517
rect 4305 -1551 4339 -1517
rect 4373 -1534 4492 -1517
rect 4526 -1534 4670 -1500
rect 4704 -1517 5312 -1500
rect 4704 -1534 4823 -1517
rect 4373 -1551 4823 -1534
rect 4857 -1551 4891 -1517
rect 4925 -1551 5091 -1517
rect 5125 -1551 5159 -1517
rect 5193 -1534 5312 -1517
rect 5346 -1534 5490 -1500
rect 5524 -1517 6132 -1500
rect 5524 -1534 5643 -1517
rect 5193 -1551 5643 -1534
rect 5677 -1551 5711 -1517
rect 5745 -1551 5911 -1517
rect 5945 -1551 5979 -1517
rect 6013 -1534 6132 -1517
rect 6166 -1534 6310 -1500
rect 6344 -1517 6952 -1500
rect 6344 -1534 6463 -1517
rect 6013 -1551 6463 -1534
rect 6497 -1551 6531 -1517
rect 6565 -1551 6731 -1517
rect 6765 -1551 6799 -1517
rect 6833 -1534 6952 -1517
rect 6986 -1534 8620 -1500
rect 6833 -1551 8620 -1534
rect -1110 -1568 8620 -1551
rect -1110 -1570 -1070 -1568
rect -1104 -1602 -1070 -1570
rect -1036 -1570 -428 -1568
rect -1036 -1602 -1003 -1570
rect -1104 -1802 -1003 -1602
rect -1104 -1830 -1070 -1802
rect -1110 -1836 -1070 -1830
rect -1036 -1830 -1003 -1802
rect -941 -1585 -869 -1570
rect -941 -1619 -917 -1585
rect -883 -1619 -869 -1585
rect -941 -1785 -869 -1619
rect -595 -1585 -523 -1570
rect -595 -1619 -581 -1585
rect -547 -1619 -523 -1585
rect -811 -1637 -653 -1623
rect -811 -1671 -797 -1637
rect -763 -1651 -701 -1637
rect -667 -1671 -653 -1637
rect -811 -1733 -783 -1671
rect -681 -1733 -653 -1671
rect -811 -1767 -797 -1733
rect -763 -1767 -701 -1753
rect -667 -1767 -653 -1733
rect -811 -1781 -653 -1767
rect -941 -1819 -917 -1785
rect -883 -1819 -869 -1785
rect -941 -1830 -869 -1819
rect -595 -1785 -523 -1619
rect -595 -1819 -581 -1785
rect -547 -1819 -523 -1785
rect -595 -1830 -523 -1819
rect -461 -1602 -428 -1570
rect -394 -1570 -250 -1568
rect -394 -1602 -360 -1570
rect -461 -1802 -360 -1602
rect -461 -1830 -428 -1802
rect -1036 -1836 -428 -1830
rect -394 -1830 -360 -1802
rect -284 -1602 -250 -1570
rect -216 -1570 392 -1568
rect -216 -1602 -183 -1570
rect -284 -1802 -183 -1602
rect -284 -1830 -250 -1802
rect -394 -1836 -250 -1830
rect -216 -1830 -183 -1802
rect -121 -1585 -49 -1570
rect -121 -1619 -97 -1585
rect -63 -1619 -49 -1585
rect -121 -1785 -49 -1619
rect 225 -1585 297 -1570
rect 225 -1619 239 -1585
rect 273 -1619 297 -1585
rect 9 -1637 167 -1623
rect 9 -1671 23 -1637
rect 57 -1651 119 -1637
rect 153 -1671 167 -1637
rect 9 -1733 37 -1671
rect 139 -1733 167 -1671
rect 9 -1767 23 -1733
rect 57 -1767 119 -1753
rect 153 -1767 167 -1733
rect 9 -1781 167 -1767
rect -121 -1819 -97 -1785
rect -63 -1819 -49 -1785
rect -121 -1830 -49 -1819
rect 225 -1785 297 -1619
rect 225 -1819 239 -1785
rect 273 -1819 297 -1785
rect 225 -1830 297 -1819
rect 359 -1602 392 -1570
rect 426 -1570 570 -1568
rect 426 -1602 460 -1570
rect 359 -1802 460 -1602
rect 359 -1830 392 -1802
rect -216 -1836 392 -1830
rect 426 -1830 460 -1802
rect 536 -1602 570 -1570
rect 604 -1570 1212 -1568
rect 604 -1602 637 -1570
rect 536 -1802 637 -1602
rect 536 -1830 570 -1802
rect 426 -1836 570 -1830
rect 604 -1830 637 -1802
rect 699 -1585 771 -1570
rect 699 -1619 723 -1585
rect 757 -1619 771 -1585
rect 699 -1785 771 -1619
rect 1045 -1585 1117 -1570
rect 1045 -1619 1059 -1585
rect 1093 -1619 1117 -1585
rect 829 -1637 987 -1623
rect 829 -1671 843 -1637
rect 877 -1651 939 -1637
rect 973 -1671 987 -1637
rect 829 -1733 857 -1671
rect 959 -1733 987 -1671
rect 829 -1767 843 -1733
rect 877 -1767 939 -1753
rect 973 -1767 987 -1733
rect 829 -1781 987 -1767
rect 699 -1819 723 -1785
rect 757 -1819 771 -1785
rect 699 -1830 771 -1819
rect 1045 -1785 1117 -1619
rect 1045 -1819 1059 -1785
rect 1093 -1819 1117 -1785
rect 1045 -1830 1117 -1819
rect 1179 -1602 1212 -1570
rect 1246 -1570 1390 -1568
rect 1246 -1602 1280 -1570
rect 1179 -1802 1280 -1602
rect 1179 -1830 1212 -1802
rect 604 -1836 1212 -1830
rect 1246 -1830 1280 -1802
rect 1356 -1602 1390 -1570
rect 1424 -1570 2032 -1568
rect 1424 -1602 1457 -1570
rect 1356 -1802 1457 -1602
rect 1356 -1830 1390 -1802
rect 1246 -1836 1390 -1830
rect 1424 -1830 1457 -1802
rect 1519 -1585 1591 -1570
rect 1519 -1619 1543 -1585
rect 1577 -1619 1591 -1585
rect 1519 -1785 1591 -1619
rect 1865 -1585 1937 -1570
rect 1865 -1619 1879 -1585
rect 1913 -1619 1937 -1585
rect 1649 -1637 1807 -1623
rect 1649 -1671 1663 -1637
rect 1697 -1651 1759 -1637
rect 1793 -1671 1807 -1637
rect 1649 -1733 1677 -1671
rect 1779 -1733 1807 -1671
rect 1649 -1767 1663 -1733
rect 1697 -1767 1759 -1753
rect 1793 -1767 1807 -1733
rect 1649 -1781 1807 -1767
rect 1519 -1819 1543 -1785
rect 1577 -1819 1591 -1785
rect 1519 -1830 1591 -1819
rect 1865 -1785 1937 -1619
rect 1865 -1819 1879 -1785
rect 1913 -1819 1937 -1785
rect 1865 -1830 1937 -1819
rect 1999 -1602 2032 -1570
rect 2066 -1570 2210 -1568
rect 2066 -1602 2100 -1570
rect 1999 -1802 2100 -1602
rect 1999 -1830 2032 -1802
rect 1424 -1836 2032 -1830
rect 2066 -1830 2100 -1802
rect 2176 -1602 2210 -1570
rect 2244 -1570 2852 -1568
rect 2244 -1602 2277 -1570
rect 2176 -1802 2277 -1602
rect 2176 -1830 2210 -1802
rect 2066 -1836 2210 -1830
rect 2244 -1830 2277 -1802
rect 2339 -1585 2411 -1570
rect 2339 -1619 2363 -1585
rect 2397 -1619 2411 -1585
rect 2339 -1785 2411 -1619
rect 2685 -1585 2757 -1570
rect 2685 -1619 2699 -1585
rect 2733 -1619 2757 -1585
rect 2469 -1637 2627 -1623
rect 2469 -1671 2483 -1637
rect 2517 -1651 2579 -1637
rect 2613 -1671 2627 -1637
rect 2469 -1733 2497 -1671
rect 2599 -1733 2627 -1671
rect 2469 -1767 2483 -1733
rect 2517 -1767 2579 -1753
rect 2613 -1767 2627 -1733
rect 2469 -1781 2627 -1767
rect 2339 -1819 2363 -1785
rect 2397 -1819 2411 -1785
rect 2339 -1830 2411 -1819
rect 2685 -1785 2757 -1619
rect 2685 -1819 2699 -1785
rect 2733 -1819 2757 -1785
rect 2685 -1830 2757 -1819
rect 2819 -1602 2852 -1570
rect 2886 -1570 3030 -1568
rect 2886 -1602 2920 -1570
rect 2819 -1802 2920 -1602
rect 2819 -1830 2852 -1802
rect 2244 -1836 2852 -1830
rect 2886 -1830 2920 -1802
rect 2996 -1602 3030 -1570
rect 3064 -1570 3672 -1568
rect 3064 -1602 3097 -1570
rect 2996 -1802 3097 -1602
rect 2996 -1830 3030 -1802
rect 2886 -1836 3030 -1830
rect 3064 -1830 3097 -1802
rect 3159 -1585 3231 -1570
rect 3159 -1619 3183 -1585
rect 3217 -1619 3231 -1585
rect 3159 -1785 3231 -1619
rect 3505 -1585 3577 -1570
rect 3505 -1619 3519 -1585
rect 3553 -1619 3577 -1585
rect 3289 -1637 3447 -1623
rect 3289 -1671 3303 -1637
rect 3337 -1651 3399 -1637
rect 3433 -1671 3447 -1637
rect 3289 -1733 3317 -1671
rect 3419 -1733 3447 -1671
rect 3289 -1767 3303 -1733
rect 3337 -1767 3399 -1753
rect 3433 -1767 3447 -1733
rect 3289 -1781 3447 -1767
rect 3159 -1819 3183 -1785
rect 3217 -1819 3231 -1785
rect 3159 -1830 3231 -1819
rect 3505 -1785 3577 -1619
rect 3505 -1819 3519 -1785
rect 3553 -1819 3577 -1785
rect 3505 -1830 3577 -1819
rect 3639 -1602 3672 -1570
rect 3706 -1570 3850 -1568
rect 3706 -1602 3740 -1570
rect 3639 -1802 3740 -1602
rect 3639 -1830 3672 -1802
rect 3064 -1836 3672 -1830
rect 3706 -1830 3740 -1802
rect 3816 -1602 3850 -1570
rect 3884 -1570 4492 -1568
rect 3884 -1602 3917 -1570
rect 3816 -1802 3917 -1602
rect 3816 -1830 3850 -1802
rect 3706 -1836 3850 -1830
rect 3884 -1830 3917 -1802
rect 3979 -1585 4051 -1570
rect 3979 -1619 4003 -1585
rect 4037 -1619 4051 -1585
rect 3979 -1785 4051 -1619
rect 4325 -1585 4397 -1570
rect 4325 -1619 4339 -1585
rect 4373 -1619 4397 -1585
rect 4109 -1637 4267 -1623
rect 4109 -1671 4123 -1637
rect 4157 -1651 4219 -1637
rect 4253 -1671 4267 -1637
rect 4109 -1733 4137 -1671
rect 4239 -1733 4267 -1671
rect 4109 -1767 4123 -1733
rect 4157 -1767 4219 -1753
rect 4253 -1767 4267 -1733
rect 4109 -1781 4267 -1767
rect 3979 -1819 4003 -1785
rect 4037 -1819 4051 -1785
rect 3979 -1830 4051 -1819
rect 4325 -1785 4397 -1619
rect 4325 -1819 4339 -1785
rect 4373 -1819 4397 -1785
rect 4325 -1830 4397 -1819
rect 4459 -1602 4492 -1570
rect 4526 -1570 4670 -1568
rect 4526 -1602 4560 -1570
rect 4459 -1802 4560 -1602
rect 4459 -1830 4492 -1802
rect 3884 -1836 4492 -1830
rect 4526 -1830 4560 -1802
rect 4636 -1602 4670 -1570
rect 4704 -1570 5312 -1568
rect 4704 -1602 4737 -1570
rect 4636 -1802 4737 -1602
rect 4636 -1830 4670 -1802
rect 4526 -1836 4670 -1830
rect 4704 -1830 4737 -1802
rect 4799 -1585 4871 -1570
rect 4799 -1619 4823 -1585
rect 4857 -1619 4871 -1585
rect 4799 -1785 4871 -1619
rect 5145 -1585 5217 -1570
rect 5145 -1619 5159 -1585
rect 5193 -1619 5217 -1585
rect 4929 -1637 5087 -1623
rect 4929 -1671 4943 -1637
rect 4977 -1651 5039 -1637
rect 5073 -1671 5087 -1637
rect 4929 -1733 4957 -1671
rect 5059 -1733 5087 -1671
rect 4929 -1767 4943 -1733
rect 4977 -1767 5039 -1753
rect 5073 -1767 5087 -1733
rect 4929 -1781 5087 -1767
rect 4799 -1819 4823 -1785
rect 4857 -1819 4871 -1785
rect 4799 -1830 4871 -1819
rect 5145 -1785 5217 -1619
rect 5145 -1819 5159 -1785
rect 5193 -1819 5217 -1785
rect 5145 -1830 5217 -1819
rect 5279 -1602 5312 -1570
rect 5346 -1570 5490 -1568
rect 5346 -1602 5380 -1570
rect 5279 -1802 5380 -1602
rect 5279 -1830 5312 -1802
rect 4704 -1836 5312 -1830
rect 5346 -1830 5380 -1802
rect 5456 -1602 5490 -1570
rect 5524 -1570 6132 -1568
rect 5524 -1602 5557 -1570
rect 5456 -1802 5557 -1602
rect 5456 -1830 5490 -1802
rect 5346 -1836 5490 -1830
rect 5524 -1830 5557 -1802
rect 5619 -1585 5691 -1570
rect 5619 -1619 5643 -1585
rect 5677 -1619 5691 -1585
rect 5619 -1785 5691 -1619
rect 5965 -1585 6037 -1570
rect 5965 -1619 5979 -1585
rect 6013 -1619 6037 -1585
rect 5749 -1637 5907 -1623
rect 5749 -1671 5763 -1637
rect 5797 -1651 5859 -1637
rect 5893 -1671 5907 -1637
rect 5749 -1733 5777 -1671
rect 5879 -1733 5907 -1671
rect 5749 -1767 5763 -1733
rect 5797 -1767 5859 -1753
rect 5893 -1767 5907 -1733
rect 5749 -1781 5907 -1767
rect 5619 -1819 5643 -1785
rect 5677 -1819 5691 -1785
rect 5619 -1830 5691 -1819
rect 5965 -1785 6037 -1619
rect 5965 -1819 5979 -1785
rect 6013 -1819 6037 -1785
rect 5965 -1830 6037 -1819
rect 6099 -1602 6132 -1570
rect 6166 -1570 6310 -1568
rect 6166 -1602 6200 -1570
rect 6099 -1802 6200 -1602
rect 6099 -1830 6132 -1802
rect 5524 -1836 6132 -1830
rect 6166 -1830 6200 -1802
rect 6276 -1602 6310 -1570
rect 6344 -1570 6952 -1568
rect 6344 -1602 6377 -1570
rect 6276 -1802 6377 -1602
rect 6276 -1830 6310 -1802
rect 6166 -1836 6310 -1830
rect 6344 -1830 6377 -1802
rect 6439 -1585 6511 -1570
rect 6439 -1619 6463 -1585
rect 6497 -1619 6511 -1585
rect 6439 -1785 6511 -1619
rect 6785 -1585 6857 -1570
rect 6785 -1619 6799 -1585
rect 6833 -1619 6857 -1585
rect 6569 -1637 6727 -1623
rect 6569 -1671 6583 -1637
rect 6617 -1651 6679 -1637
rect 6713 -1671 6727 -1637
rect 6569 -1733 6597 -1671
rect 6699 -1733 6727 -1671
rect 6569 -1767 6583 -1733
rect 6617 -1767 6679 -1753
rect 6713 -1767 6727 -1733
rect 6569 -1781 6727 -1767
rect 6439 -1819 6463 -1785
rect 6497 -1819 6511 -1785
rect 6439 -1830 6511 -1819
rect 6785 -1785 6857 -1619
rect 6785 -1819 6799 -1785
rect 6833 -1819 6857 -1785
rect 6785 -1830 6857 -1819
rect 6919 -1602 6952 -1570
rect 6986 -1602 8620 -1568
rect 6919 -1630 8620 -1602
rect 8760 -1630 8790 -1170
rect 16330 -1340 16580 -900
rect 6919 -1660 8790 -1630
rect 6919 -1802 7020 -1660
rect 6919 -1830 6952 -1802
rect 6344 -1836 6952 -1830
rect 6986 -1830 7020 -1802
rect 6986 -1836 7030 -1830
rect -1110 -1853 7030 -1836
rect -1110 -1870 -917 -1853
rect -1110 -1904 -1070 -1870
rect -1036 -1887 -917 -1870
rect -883 -1887 -849 -1853
rect -815 -1887 -649 -1853
rect -615 -1887 -581 -1853
rect -547 -1870 -97 -1853
rect -547 -1887 -428 -1870
rect -1036 -1904 -428 -1887
rect -394 -1904 -250 -1870
rect -216 -1887 -97 -1870
rect -63 -1887 -29 -1853
rect 5 -1887 171 -1853
rect 205 -1887 239 -1853
rect 273 -1870 723 -1853
rect 273 -1887 392 -1870
rect -216 -1904 392 -1887
rect 426 -1904 570 -1870
rect 604 -1887 723 -1870
rect 757 -1887 791 -1853
rect 825 -1887 991 -1853
rect 1025 -1887 1059 -1853
rect 1093 -1870 1543 -1853
rect 1093 -1887 1212 -1870
rect 604 -1904 1212 -1887
rect 1246 -1904 1390 -1870
rect 1424 -1887 1543 -1870
rect 1577 -1887 1611 -1853
rect 1645 -1887 1811 -1853
rect 1845 -1887 1879 -1853
rect 1913 -1870 2363 -1853
rect 1913 -1887 2032 -1870
rect 1424 -1904 2032 -1887
rect 2066 -1904 2210 -1870
rect 2244 -1887 2363 -1870
rect 2397 -1887 2431 -1853
rect 2465 -1887 2631 -1853
rect 2665 -1887 2699 -1853
rect 2733 -1870 3183 -1853
rect 2733 -1887 2852 -1870
rect 2244 -1904 2852 -1887
rect 2886 -1904 3030 -1870
rect 3064 -1887 3183 -1870
rect 3217 -1887 3251 -1853
rect 3285 -1887 3451 -1853
rect 3485 -1887 3519 -1853
rect 3553 -1870 4003 -1853
rect 3553 -1887 3672 -1870
rect 3064 -1904 3672 -1887
rect 3706 -1904 3850 -1870
rect 3884 -1887 4003 -1870
rect 4037 -1887 4071 -1853
rect 4105 -1887 4271 -1853
rect 4305 -1887 4339 -1853
rect 4373 -1870 4823 -1853
rect 4373 -1887 4492 -1870
rect 3884 -1904 4492 -1887
rect 4526 -1904 4670 -1870
rect 4704 -1887 4823 -1870
rect 4857 -1887 4891 -1853
rect 4925 -1887 5091 -1853
rect 5125 -1887 5159 -1853
rect 5193 -1870 5643 -1853
rect 5193 -1887 5312 -1870
rect 4704 -1904 5312 -1887
rect 5346 -1904 5490 -1870
rect 5524 -1887 5643 -1870
rect 5677 -1887 5711 -1853
rect 5745 -1887 5911 -1853
rect 5945 -1887 5979 -1853
rect 6013 -1870 6463 -1853
rect 6013 -1887 6132 -1870
rect 5524 -1904 6132 -1887
rect 6166 -1904 6310 -1870
rect 6344 -1887 6463 -1870
rect 6497 -1887 6531 -1853
rect 6565 -1887 6731 -1853
rect 6765 -1887 6799 -1853
rect 6833 -1870 7030 -1853
rect 6833 -1887 6952 -1870
rect 6344 -1904 6952 -1887
rect 6986 -1904 7030 -1870
rect -1110 -1938 7030 -1904
rect -1110 -1972 -1070 -1938
rect -1036 -1972 -428 -1938
rect -394 -1972 -250 -1938
rect -216 -1972 392 -1938
rect 426 -1972 570 -1938
rect 604 -1972 1212 -1938
rect 1246 -1972 1390 -1938
rect 1424 -1972 2032 -1938
rect 2066 -1972 2210 -1938
rect 2244 -1972 2852 -1938
rect 2886 -1972 3030 -1938
rect 3064 -1972 3672 -1938
rect 3706 -1972 3850 -1938
rect 3884 -1972 4492 -1938
rect 4526 -1972 4670 -1938
rect 4704 -1972 5312 -1938
rect 5346 -1972 5490 -1938
rect 5524 -1972 6132 -1938
rect 6166 -1972 6310 -1938
rect 6344 -1972 6952 -1938
rect 6986 -1972 7030 -1938
rect -1110 -2006 7030 -1972
rect -1110 -2040 -1070 -2006
rect -1036 -2040 -1002 -2006
rect -968 -2040 -934 -2006
rect -900 -2040 -866 -2006
rect -832 -2040 -632 -2006
rect -598 -2040 -564 -2006
rect -530 -2040 -496 -2006
rect -462 -2040 -428 -2006
rect -394 -2040 -250 -2006
rect -216 -2040 -182 -2006
rect -148 -2040 -114 -2006
rect -80 -2040 -46 -2006
rect -12 -2040 188 -2006
rect 222 -2040 256 -2006
rect 290 -2040 324 -2006
rect 358 -2040 392 -2006
rect 426 -2040 570 -2006
rect 604 -2040 638 -2006
rect 672 -2040 706 -2006
rect 740 -2040 774 -2006
rect 808 -2040 1008 -2006
rect 1042 -2040 1076 -2006
rect 1110 -2040 1144 -2006
rect 1178 -2040 1212 -2006
rect 1246 -2040 1390 -2006
rect 1424 -2040 1458 -2006
rect 1492 -2040 1526 -2006
rect 1560 -2040 1594 -2006
rect 1628 -2040 1828 -2006
rect 1862 -2040 1896 -2006
rect 1930 -2040 1964 -2006
rect 1998 -2040 2032 -2006
rect 2066 -2040 2210 -2006
rect 2244 -2040 2278 -2006
rect 2312 -2040 2346 -2006
rect 2380 -2040 2414 -2006
rect 2448 -2040 2648 -2006
rect 2682 -2040 2716 -2006
rect 2750 -2040 2784 -2006
rect 2818 -2040 2852 -2006
rect 2886 -2040 3030 -2006
rect 3064 -2040 3098 -2006
rect 3132 -2040 3166 -2006
rect 3200 -2040 3234 -2006
rect 3268 -2040 3468 -2006
rect 3502 -2040 3536 -2006
rect 3570 -2040 3604 -2006
rect 3638 -2040 3672 -2006
rect 3706 -2040 3850 -2006
rect 3884 -2040 3918 -2006
rect 3952 -2040 3986 -2006
rect 4020 -2040 4054 -2006
rect 4088 -2040 4288 -2006
rect 4322 -2040 4356 -2006
rect 4390 -2040 4424 -2006
rect 4458 -2040 4492 -2006
rect 4526 -2040 4670 -2006
rect 4704 -2040 4738 -2006
rect 4772 -2040 4806 -2006
rect 4840 -2040 4874 -2006
rect 4908 -2040 5108 -2006
rect 5142 -2040 5176 -2006
rect 5210 -2040 5244 -2006
rect 5278 -2040 5312 -2006
rect 5346 -2040 5490 -2006
rect 5524 -2040 5558 -2006
rect 5592 -2040 5626 -2006
rect 5660 -2040 5694 -2006
rect 5728 -2040 5928 -2006
rect 5962 -2040 5996 -2006
rect 6030 -2040 6064 -2006
rect 6098 -2040 6132 -2006
rect 6166 -2040 6310 -2006
rect 6344 -2040 6378 -2006
rect 6412 -2040 6446 -2006
rect 6480 -2040 6514 -2006
rect 6548 -2040 6748 -2006
rect 6782 -2040 6816 -2006
rect 6850 -2040 6884 -2006
rect 6918 -2040 6952 -2006
rect 6986 -2040 7030 -2006
rect -1110 -2184 7030 -2040
rect -1110 -2218 -1070 -2184
rect -1036 -2218 -1002 -2184
rect -968 -2218 -934 -2184
rect -900 -2218 -866 -2184
rect -832 -2218 -632 -2184
rect -598 -2218 -564 -2184
rect -530 -2218 -496 -2184
rect -462 -2218 -428 -2184
rect -394 -2218 -250 -2184
rect -216 -2218 -182 -2184
rect -148 -2218 -114 -2184
rect -80 -2218 -46 -2184
rect -12 -2218 188 -2184
rect 222 -2218 256 -2184
rect 290 -2218 324 -2184
rect 358 -2218 392 -2184
rect 426 -2218 570 -2184
rect 604 -2218 638 -2184
rect 672 -2218 706 -2184
rect 740 -2218 774 -2184
rect 808 -2218 1008 -2184
rect 1042 -2218 1076 -2184
rect 1110 -2218 1144 -2184
rect 1178 -2218 1212 -2184
rect 1246 -2218 1390 -2184
rect 1424 -2218 1458 -2184
rect 1492 -2218 1526 -2184
rect 1560 -2218 1594 -2184
rect 1628 -2218 1828 -2184
rect 1862 -2218 1896 -2184
rect 1930 -2218 1964 -2184
rect 1998 -2218 2032 -2184
rect 2066 -2218 2210 -2184
rect 2244 -2218 2278 -2184
rect 2312 -2218 2346 -2184
rect 2380 -2218 2414 -2184
rect 2448 -2218 2648 -2184
rect 2682 -2218 2716 -2184
rect 2750 -2218 2784 -2184
rect 2818 -2218 2852 -2184
rect 2886 -2218 3030 -2184
rect 3064 -2218 3098 -2184
rect 3132 -2218 3166 -2184
rect 3200 -2218 3234 -2184
rect 3268 -2218 3468 -2184
rect 3502 -2218 3536 -2184
rect 3570 -2218 3604 -2184
rect 3638 -2218 3672 -2184
rect 3706 -2218 3850 -2184
rect 3884 -2218 3918 -2184
rect 3952 -2218 3986 -2184
rect 4020 -2218 4054 -2184
rect 4088 -2218 4288 -2184
rect 4322 -2218 4356 -2184
rect 4390 -2218 4424 -2184
rect 4458 -2218 4492 -2184
rect 4526 -2218 4670 -2184
rect 4704 -2218 4738 -2184
rect 4772 -2218 4806 -2184
rect 4840 -2218 4874 -2184
rect 4908 -2218 5108 -2184
rect 5142 -2218 5176 -2184
rect 5210 -2218 5244 -2184
rect 5278 -2218 5312 -2184
rect 5346 -2218 5490 -2184
rect 5524 -2218 5558 -2184
rect 5592 -2218 5626 -2184
rect 5660 -2218 5694 -2184
rect 5728 -2218 5928 -2184
rect 5962 -2218 5996 -2184
rect 6030 -2218 6064 -2184
rect 6098 -2218 6132 -2184
rect 6166 -2218 6310 -2184
rect 6344 -2218 6378 -2184
rect 6412 -2218 6446 -2184
rect 6480 -2218 6514 -2184
rect 6548 -2218 6748 -2184
rect 6782 -2218 6816 -2184
rect 6850 -2218 6884 -2184
rect 6918 -2218 6952 -2184
rect 6986 -2218 7030 -2184
rect -1110 -2252 7030 -2218
rect -1110 -2286 -1070 -2252
rect -1036 -2286 -428 -2252
rect -394 -2286 -250 -2252
rect -216 -2286 392 -2252
rect 426 -2286 570 -2252
rect 604 -2286 1212 -2252
rect 1246 -2286 1390 -2252
rect 1424 -2286 2032 -2252
rect 2066 -2286 2210 -2252
rect 2244 -2286 2852 -2252
rect 2886 -2286 3030 -2252
rect 3064 -2286 3672 -2252
rect 3706 -2286 3850 -2252
rect 3884 -2286 4492 -2252
rect 4526 -2286 4670 -2252
rect 4704 -2286 5312 -2252
rect 5346 -2286 5490 -2252
rect 5524 -2286 6132 -2252
rect 6166 -2286 6310 -2252
rect 6344 -2286 6952 -2252
rect 6986 -2286 7030 -2252
rect -1110 -2320 7030 -2286
rect -1110 -2354 -1070 -2320
rect -1036 -2337 -428 -2320
rect -1036 -2354 -917 -2337
rect -1110 -2371 -917 -2354
rect -883 -2371 -849 -2337
rect -815 -2371 -649 -2337
rect -615 -2371 -581 -2337
rect -547 -2354 -428 -2337
rect -394 -2354 -250 -2320
rect -216 -2337 392 -2320
rect -216 -2354 -97 -2337
rect -547 -2371 -97 -2354
rect -63 -2371 -29 -2337
rect 5 -2371 171 -2337
rect 205 -2371 239 -2337
rect 273 -2354 392 -2337
rect 426 -2354 570 -2320
rect 604 -2337 1212 -2320
rect 604 -2354 723 -2337
rect 273 -2371 723 -2354
rect 757 -2371 791 -2337
rect 825 -2371 991 -2337
rect 1025 -2371 1059 -2337
rect 1093 -2354 1212 -2337
rect 1246 -2354 1390 -2320
rect 1424 -2337 2032 -2320
rect 1424 -2354 1543 -2337
rect 1093 -2371 1543 -2354
rect 1577 -2371 1611 -2337
rect 1645 -2371 1811 -2337
rect 1845 -2371 1879 -2337
rect 1913 -2354 2032 -2337
rect 2066 -2354 2210 -2320
rect 2244 -2337 2852 -2320
rect 2244 -2354 2363 -2337
rect 1913 -2371 2363 -2354
rect 2397 -2371 2431 -2337
rect 2465 -2371 2631 -2337
rect 2665 -2371 2699 -2337
rect 2733 -2354 2852 -2337
rect 2886 -2354 3030 -2320
rect 3064 -2337 3672 -2320
rect 3064 -2354 3183 -2337
rect 2733 -2371 3183 -2354
rect 3217 -2371 3251 -2337
rect 3285 -2371 3451 -2337
rect 3485 -2371 3519 -2337
rect 3553 -2354 3672 -2337
rect 3706 -2354 3850 -2320
rect 3884 -2337 4492 -2320
rect 3884 -2354 4003 -2337
rect 3553 -2371 4003 -2354
rect 4037 -2371 4071 -2337
rect 4105 -2371 4271 -2337
rect 4305 -2371 4339 -2337
rect 4373 -2354 4492 -2337
rect 4526 -2354 4670 -2320
rect 4704 -2337 5312 -2320
rect 4704 -2354 4823 -2337
rect 4373 -2371 4823 -2354
rect 4857 -2371 4891 -2337
rect 4925 -2371 5091 -2337
rect 5125 -2371 5159 -2337
rect 5193 -2354 5312 -2337
rect 5346 -2354 5490 -2320
rect 5524 -2337 6132 -2320
rect 5524 -2354 5643 -2337
rect 5193 -2371 5643 -2354
rect 5677 -2371 5711 -2337
rect 5745 -2371 5911 -2337
rect 5945 -2371 5979 -2337
rect 6013 -2354 6132 -2337
rect 6166 -2354 6310 -2320
rect 6344 -2337 6952 -2320
rect 6344 -2354 6463 -2337
rect 6013 -2371 6463 -2354
rect 6497 -2371 6531 -2337
rect 6565 -2371 6731 -2337
rect 6765 -2371 6799 -2337
rect 6833 -2354 6952 -2337
rect 6986 -2354 7030 -2320
rect 6833 -2371 7030 -2354
rect -1110 -2388 7030 -2371
rect -1110 -2390 -1070 -2388
rect -1104 -2422 -1070 -2390
rect -1036 -2390 -428 -2388
rect -1036 -2422 -1003 -2390
rect -1104 -2622 -1003 -2422
rect -1104 -2650 -1070 -2622
rect -1110 -2656 -1070 -2650
rect -1036 -2650 -1003 -2622
rect -941 -2405 -869 -2390
rect -941 -2439 -917 -2405
rect -883 -2439 -869 -2405
rect -941 -2605 -869 -2439
rect -595 -2405 -523 -2390
rect -595 -2439 -581 -2405
rect -547 -2439 -523 -2405
rect -811 -2457 -653 -2443
rect -811 -2491 -797 -2457
rect -763 -2471 -701 -2457
rect -667 -2491 -653 -2457
rect -811 -2553 -783 -2491
rect -681 -2553 -653 -2491
rect -811 -2587 -797 -2553
rect -763 -2587 -701 -2573
rect -667 -2587 -653 -2553
rect -811 -2601 -653 -2587
rect -941 -2639 -917 -2605
rect -883 -2639 -869 -2605
rect -941 -2650 -869 -2639
rect -595 -2605 -523 -2439
rect -595 -2639 -581 -2605
rect -547 -2639 -523 -2605
rect -595 -2650 -523 -2639
rect -461 -2422 -428 -2390
rect -394 -2390 -250 -2388
rect -394 -2422 -360 -2390
rect -461 -2622 -360 -2422
rect -461 -2650 -428 -2622
rect -1036 -2656 -428 -2650
rect -394 -2650 -360 -2622
rect -284 -2422 -250 -2390
rect -216 -2390 392 -2388
rect -216 -2422 -183 -2390
rect -284 -2622 -183 -2422
rect -284 -2650 -250 -2622
rect -394 -2656 -250 -2650
rect -216 -2650 -183 -2622
rect -121 -2405 -49 -2390
rect -121 -2439 -97 -2405
rect -63 -2439 -49 -2405
rect -121 -2605 -49 -2439
rect 225 -2405 297 -2390
rect 225 -2439 239 -2405
rect 273 -2439 297 -2405
rect 9 -2457 167 -2443
rect 9 -2491 23 -2457
rect 57 -2471 119 -2457
rect 153 -2491 167 -2457
rect 9 -2553 37 -2491
rect 139 -2553 167 -2491
rect 9 -2587 23 -2553
rect 57 -2587 119 -2573
rect 153 -2587 167 -2553
rect 9 -2601 167 -2587
rect -121 -2639 -97 -2605
rect -63 -2639 -49 -2605
rect -121 -2650 -49 -2639
rect 225 -2605 297 -2439
rect 225 -2639 239 -2605
rect 273 -2639 297 -2605
rect 225 -2650 297 -2639
rect 359 -2422 392 -2390
rect 426 -2390 570 -2388
rect 426 -2422 460 -2390
rect 359 -2622 460 -2422
rect 359 -2650 392 -2622
rect -216 -2656 392 -2650
rect 426 -2650 460 -2622
rect 536 -2422 570 -2390
rect 604 -2390 1212 -2388
rect 604 -2422 637 -2390
rect 536 -2622 637 -2422
rect 536 -2650 570 -2622
rect 426 -2656 570 -2650
rect 604 -2650 637 -2622
rect 699 -2405 771 -2390
rect 699 -2439 723 -2405
rect 757 -2439 771 -2405
rect 699 -2605 771 -2439
rect 1045 -2405 1117 -2390
rect 1045 -2439 1059 -2405
rect 1093 -2439 1117 -2405
rect 829 -2457 987 -2443
rect 829 -2491 843 -2457
rect 877 -2471 939 -2457
rect 973 -2491 987 -2457
rect 829 -2553 857 -2491
rect 959 -2553 987 -2491
rect 829 -2587 843 -2553
rect 877 -2587 939 -2573
rect 973 -2587 987 -2553
rect 829 -2601 987 -2587
rect 699 -2639 723 -2605
rect 757 -2639 771 -2605
rect 699 -2650 771 -2639
rect 1045 -2605 1117 -2439
rect 1045 -2639 1059 -2605
rect 1093 -2639 1117 -2605
rect 1045 -2650 1117 -2639
rect 1179 -2422 1212 -2390
rect 1246 -2390 1390 -2388
rect 1246 -2422 1280 -2390
rect 1179 -2622 1280 -2422
rect 1179 -2650 1212 -2622
rect 604 -2656 1212 -2650
rect 1246 -2650 1280 -2622
rect 1356 -2422 1390 -2390
rect 1424 -2390 2032 -2388
rect 1424 -2422 1457 -2390
rect 1356 -2622 1457 -2422
rect 1356 -2650 1390 -2622
rect 1246 -2656 1390 -2650
rect 1424 -2650 1457 -2622
rect 1519 -2405 1591 -2390
rect 1519 -2439 1543 -2405
rect 1577 -2439 1591 -2405
rect 1519 -2605 1591 -2439
rect 1865 -2405 1937 -2390
rect 1865 -2439 1879 -2405
rect 1913 -2439 1937 -2405
rect 1649 -2457 1807 -2443
rect 1649 -2491 1663 -2457
rect 1697 -2471 1759 -2457
rect 1793 -2491 1807 -2457
rect 1649 -2553 1677 -2491
rect 1779 -2553 1807 -2491
rect 1649 -2587 1663 -2553
rect 1697 -2587 1759 -2573
rect 1793 -2587 1807 -2553
rect 1649 -2601 1807 -2587
rect 1519 -2639 1543 -2605
rect 1577 -2639 1591 -2605
rect 1519 -2650 1591 -2639
rect 1865 -2605 1937 -2439
rect 1865 -2639 1879 -2605
rect 1913 -2639 1937 -2605
rect 1865 -2650 1937 -2639
rect 1999 -2422 2032 -2390
rect 2066 -2390 2210 -2388
rect 2066 -2422 2100 -2390
rect 1999 -2622 2100 -2422
rect 1999 -2650 2032 -2622
rect 1424 -2656 2032 -2650
rect 2066 -2650 2100 -2622
rect 2176 -2422 2210 -2390
rect 2244 -2390 2852 -2388
rect 2244 -2422 2277 -2390
rect 2176 -2622 2277 -2422
rect 2176 -2650 2210 -2622
rect 2066 -2656 2210 -2650
rect 2244 -2650 2277 -2622
rect 2339 -2405 2411 -2390
rect 2339 -2439 2363 -2405
rect 2397 -2439 2411 -2405
rect 2339 -2605 2411 -2439
rect 2685 -2405 2757 -2390
rect 2685 -2439 2699 -2405
rect 2733 -2439 2757 -2405
rect 2469 -2457 2627 -2443
rect 2469 -2491 2483 -2457
rect 2517 -2471 2579 -2457
rect 2613 -2491 2627 -2457
rect 2469 -2553 2497 -2491
rect 2599 -2553 2627 -2491
rect 2469 -2587 2483 -2553
rect 2517 -2587 2579 -2573
rect 2613 -2587 2627 -2553
rect 2469 -2601 2627 -2587
rect 2339 -2639 2363 -2605
rect 2397 -2639 2411 -2605
rect 2339 -2650 2411 -2639
rect 2685 -2605 2757 -2439
rect 2685 -2639 2699 -2605
rect 2733 -2639 2757 -2605
rect 2685 -2650 2757 -2639
rect 2819 -2422 2852 -2390
rect 2886 -2390 3030 -2388
rect 2886 -2422 2920 -2390
rect 2819 -2622 2920 -2422
rect 2819 -2650 2852 -2622
rect 2244 -2656 2852 -2650
rect 2886 -2650 2920 -2622
rect 2996 -2422 3030 -2390
rect 3064 -2390 3672 -2388
rect 3064 -2422 3097 -2390
rect 2996 -2622 3097 -2422
rect 2996 -2650 3030 -2622
rect 2886 -2656 3030 -2650
rect 3064 -2650 3097 -2622
rect 3159 -2405 3231 -2390
rect 3159 -2439 3183 -2405
rect 3217 -2439 3231 -2405
rect 3159 -2605 3231 -2439
rect 3505 -2405 3577 -2390
rect 3505 -2439 3519 -2405
rect 3553 -2439 3577 -2405
rect 3289 -2457 3447 -2443
rect 3289 -2491 3303 -2457
rect 3337 -2471 3399 -2457
rect 3433 -2491 3447 -2457
rect 3289 -2553 3317 -2491
rect 3419 -2553 3447 -2491
rect 3289 -2587 3303 -2553
rect 3337 -2587 3399 -2573
rect 3433 -2587 3447 -2553
rect 3289 -2601 3447 -2587
rect 3159 -2639 3183 -2605
rect 3217 -2639 3231 -2605
rect 3159 -2650 3231 -2639
rect 3505 -2605 3577 -2439
rect 3505 -2639 3519 -2605
rect 3553 -2639 3577 -2605
rect 3505 -2650 3577 -2639
rect 3639 -2422 3672 -2390
rect 3706 -2390 3850 -2388
rect 3706 -2422 3740 -2390
rect 3639 -2622 3740 -2422
rect 3639 -2650 3672 -2622
rect 3064 -2656 3672 -2650
rect 3706 -2650 3740 -2622
rect 3816 -2422 3850 -2390
rect 3884 -2390 4492 -2388
rect 3884 -2422 3917 -2390
rect 3816 -2622 3917 -2422
rect 3816 -2650 3850 -2622
rect 3706 -2656 3850 -2650
rect 3884 -2650 3917 -2622
rect 3979 -2405 4051 -2390
rect 3979 -2439 4003 -2405
rect 4037 -2439 4051 -2405
rect 3979 -2605 4051 -2439
rect 4325 -2405 4397 -2390
rect 4325 -2439 4339 -2405
rect 4373 -2439 4397 -2405
rect 4109 -2457 4267 -2443
rect 4109 -2491 4123 -2457
rect 4157 -2471 4219 -2457
rect 4253 -2491 4267 -2457
rect 4109 -2553 4137 -2491
rect 4239 -2553 4267 -2491
rect 4109 -2587 4123 -2553
rect 4157 -2587 4219 -2573
rect 4253 -2587 4267 -2553
rect 4109 -2601 4267 -2587
rect 3979 -2639 4003 -2605
rect 4037 -2639 4051 -2605
rect 3979 -2650 4051 -2639
rect 4325 -2605 4397 -2439
rect 4325 -2639 4339 -2605
rect 4373 -2639 4397 -2605
rect 4325 -2650 4397 -2639
rect 4459 -2422 4492 -2390
rect 4526 -2390 4670 -2388
rect 4526 -2422 4560 -2390
rect 4459 -2622 4560 -2422
rect 4459 -2650 4492 -2622
rect 3884 -2656 4492 -2650
rect 4526 -2650 4560 -2622
rect 4636 -2422 4670 -2390
rect 4704 -2390 5312 -2388
rect 4704 -2422 4737 -2390
rect 4636 -2622 4737 -2422
rect 4636 -2650 4670 -2622
rect 4526 -2656 4670 -2650
rect 4704 -2650 4737 -2622
rect 4799 -2405 4871 -2390
rect 4799 -2439 4823 -2405
rect 4857 -2439 4871 -2405
rect 4799 -2605 4871 -2439
rect 5145 -2405 5217 -2390
rect 5145 -2439 5159 -2405
rect 5193 -2439 5217 -2405
rect 4929 -2457 5087 -2443
rect 4929 -2491 4943 -2457
rect 4977 -2471 5039 -2457
rect 5073 -2491 5087 -2457
rect 4929 -2553 4957 -2491
rect 5059 -2553 5087 -2491
rect 4929 -2587 4943 -2553
rect 4977 -2587 5039 -2573
rect 5073 -2587 5087 -2553
rect 4929 -2601 5087 -2587
rect 4799 -2639 4823 -2605
rect 4857 -2639 4871 -2605
rect 4799 -2650 4871 -2639
rect 5145 -2605 5217 -2439
rect 5145 -2639 5159 -2605
rect 5193 -2639 5217 -2605
rect 5145 -2650 5217 -2639
rect 5279 -2422 5312 -2390
rect 5346 -2390 5490 -2388
rect 5346 -2422 5380 -2390
rect 5279 -2622 5380 -2422
rect 5279 -2650 5312 -2622
rect 4704 -2656 5312 -2650
rect 5346 -2650 5380 -2622
rect 5456 -2422 5490 -2390
rect 5524 -2390 6132 -2388
rect 5524 -2422 5557 -2390
rect 5456 -2622 5557 -2422
rect 5456 -2650 5490 -2622
rect 5346 -2656 5490 -2650
rect 5524 -2650 5557 -2622
rect 5619 -2405 5691 -2390
rect 5619 -2439 5643 -2405
rect 5677 -2439 5691 -2405
rect 5619 -2605 5691 -2439
rect 5965 -2405 6037 -2390
rect 5965 -2439 5979 -2405
rect 6013 -2439 6037 -2405
rect 5749 -2457 5907 -2443
rect 5749 -2491 5763 -2457
rect 5797 -2471 5859 -2457
rect 5893 -2491 5907 -2457
rect 5749 -2553 5777 -2491
rect 5879 -2553 5907 -2491
rect 5749 -2587 5763 -2553
rect 5797 -2587 5859 -2573
rect 5893 -2587 5907 -2553
rect 5749 -2601 5907 -2587
rect 5619 -2639 5643 -2605
rect 5677 -2639 5691 -2605
rect 5619 -2650 5691 -2639
rect 5965 -2605 6037 -2439
rect 5965 -2639 5979 -2605
rect 6013 -2639 6037 -2605
rect 5965 -2650 6037 -2639
rect 6099 -2422 6132 -2390
rect 6166 -2390 6310 -2388
rect 6166 -2422 6200 -2390
rect 6099 -2622 6200 -2422
rect 6099 -2650 6132 -2622
rect 5524 -2656 6132 -2650
rect 6166 -2650 6200 -2622
rect 6276 -2422 6310 -2390
rect 6344 -2390 6952 -2388
rect 6344 -2422 6377 -2390
rect 6276 -2622 6377 -2422
rect 6276 -2650 6310 -2622
rect 6166 -2656 6310 -2650
rect 6344 -2650 6377 -2622
rect 6439 -2405 6511 -2390
rect 6439 -2439 6463 -2405
rect 6497 -2439 6511 -2405
rect 6439 -2605 6511 -2439
rect 6785 -2405 6857 -2390
rect 6785 -2439 6799 -2405
rect 6833 -2439 6857 -2405
rect 6569 -2457 6727 -2443
rect 6569 -2491 6583 -2457
rect 6617 -2471 6679 -2457
rect 6713 -2491 6727 -2457
rect 6569 -2553 6597 -2491
rect 6699 -2553 6727 -2491
rect 6569 -2587 6583 -2553
rect 6617 -2587 6679 -2573
rect 6713 -2587 6727 -2553
rect 6569 -2601 6727 -2587
rect 6439 -2639 6463 -2605
rect 6497 -2639 6511 -2605
rect 6439 -2650 6511 -2639
rect 6785 -2605 6857 -2439
rect 6785 -2639 6799 -2605
rect 6833 -2639 6857 -2605
rect 6785 -2650 6857 -2639
rect 6919 -2422 6952 -2390
rect 6986 -2390 7030 -2388
rect 6986 -2422 7020 -2390
rect 6919 -2622 7020 -2422
rect 6919 -2650 6952 -2622
rect 6344 -2656 6952 -2650
rect 6986 -2650 7020 -2622
rect 6986 -2656 7030 -2650
rect -1110 -2673 7030 -2656
rect -1110 -2690 -917 -2673
rect -1110 -2724 -1070 -2690
rect -1036 -2707 -917 -2690
rect -883 -2707 -849 -2673
rect -815 -2707 -649 -2673
rect -615 -2707 -581 -2673
rect -547 -2690 -97 -2673
rect -547 -2707 -428 -2690
rect -1036 -2724 -428 -2707
rect -394 -2724 -250 -2690
rect -216 -2707 -97 -2690
rect -63 -2707 -29 -2673
rect 5 -2707 171 -2673
rect 205 -2707 239 -2673
rect 273 -2690 723 -2673
rect 273 -2707 392 -2690
rect -216 -2724 392 -2707
rect 426 -2724 570 -2690
rect 604 -2707 723 -2690
rect 757 -2707 791 -2673
rect 825 -2707 991 -2673
rect 1025 -2707 1059 -2673
rect 1093 -2690 1543 -2673
rect 1093 -2707 1212 -2690
rect 604 -2724 1212 -2707
rect 1246 -2724 1390 -2690
rect 1424 -2707 1543 -2690
rect 1577 -2707 1611 -2673
rect 1645 -2707 1811 -2673
rect 1845 -2707 1879 -2673
rect 1913 -2690 2363 -2673
rect 1913 -2707 2032 -2690
rect 1424 -2724 2032 -2707
rect 2066 -2724 2210 -2690
rect 2244 -2707 2363 -2690
rect 2397 -2707 2431 -2673
rect 2465 -2707 2631 -2673
rect 2665 -2707 2699 -2673
rect 2733 -2690 3183 -2673
rect 2733 -2707 2852 -2690
rect 2244 -2724 2852 -2707
rect 2886 -2724 3030 -2690
rect 3064 -2707 3183 -2690
rect 3217 -2707 3251 -2673
rect 3285 -2707 3451 -2673
rect 3485 -2707 3519 -2673
rect 3553 -2690 4003 -2673
rect 3553 -2707 3672 -2690
rect 3064 -2724 3672 -2707
rect 3706 -2724 3850 -2690
rect 3884 -2707 4003 -2690
rect 4037 -2707 4071 -2673
rect 4105 -2707 4271 -2673
rect 4305 -2707 4339 -2673
rect 4373 -2690 4823 -2673
rect 4373 -2707 4492 -2690
rect 3884 -2724 4492 -2707
rect 4526 -2724 4670 -2690
rect 4704 -2707 4823 -2690
rect 4857 -2707 4891 -2673
rect 4925 -2707 5091 -2673
rect 5125 -2707 5159 -2673
rect 5193 -2690 5643 -2673
rect 5193 -2707 5312 -2690
rect 4704 -2724 5312 -2707
rect 5346 -2724 5490 -2690
rect 5524 -2707 5643 -2690
rect 5677 -2707 5711 -2673
rect 5745 -2707 5911 -2673
rect 5945 -2707 5979 -2673
rect 6013 -2690 6463 -2673
rect 6013 -2707 6132 -2690
rect 5524 -2724 6132 -2707
rect 6166 -2724 6310 -2690
rect 6344 -2707 6463 -2690
rect 6497 -2707 6531 -2673
rect 6565 -2707 6731 -2673
rect 6765 -2707 6799 -2673
rect 6833 -2690 7030 -2673
rect 6833 -2707 6952 -2690
rect 6344 -2724 6952 -2707
rect 6986 -2724 7030 -2690
rect -1110 -2758 7030 -2724
rect -1110 -2792 -1070 -2758
rect -1036 -2792 -428 -2758
rect -394 -2792 -250 -2758
rect -216 -2792 392 -2758
rect 426 -2792 570 -2758
rect 604 -2792 1212 -2758
rect 1246 -2792 1390 -2758
rect 1424 -2792 2032 -2758
rect 2066 -2792 2210 -2758
rect 2244 -2792 2852 -2758
rect 2886 -2792 3030 -2758
rect 3064 -2792 3672 -2758
rect 3706 -2792 3850 -2758
rect 3884 -2792 4492 -2758
rect 4526 -2792 4670 -2758
rect 4704 -2792 5312 -2758
rect 5346 -2792 5490 -2758
rect 5524 -2792 6132 -2758
rect 6166 -2792 6310 -2758
rect 6344 -2792 6952 -2758
rect 6986 -2792 7030 -2758
rect -1110 -2826 7030 -2792
rect -1110 -2860 -1070 -2826
rect -1036 -2860 -1002 -2826
rect -968 -2860 -934 -2826
rect -900 -2860 -866 -2826
rect -832 -2860 -632 -2826
rect -598 -2860 -564 -2826
rect -530 -2860 -496 -2826
rect -462 -2860 -428 -2826
rect -394 -2860 -250 -2826
rect -216 -2860 -182 -2826
rect -148 -2860 -114 -2826
rect -80 -2860 -46 -2826
rect -12 -2860 188 -2826
rect 222 -2860 256 -2826
rect 290 -2860 324 -2826
rect 358 -2860 392 -2826
rect 426 -2860 570 -2826
rect 604 -2860 638 -2826
rect 672 -2860 706 -2826
rect 740 -2860 774 -2826
rect 808 -2860 1008 -2826
rect 1042 -2860 1076 -2826
rect 1110 -2860 1144 -2826
rect 1178 -2860 1212 -2826
rect 1246 -2860 1390 -2826
rect 1424 -2860 1458 -2826
rect 1492 -2860 1526 -2826
rect 1560 -2860 1594 -2826
rect 1628 -2860 1828 -2826
rect 1862 -2860 1896 -2826
rect 1930 -2860 1964 -2826
rect 1998 -2860 2032 -2826
rect 2066 -2860 2210 -2826
rect 2244 -2860 2278 -2826
rect 2312 -2860 2346 -2826
rect 2380 -2860 2414 -2826
rect 2448 -2860 2648 -2826
rect 2682 -2860 2716 -2826
rect 2750 -2860 2784 -2826
rect 2818 -2860 2852 -2826
rect 2886 -2860 3030 -2826
rect 3064 -2860 3098 -2826
rect 3132 -2860 3166 -2826
rect 3200 -2860 3234 -2826
rect 3268 -2860 3468 -2826
rect 3502 -2860 3536 -2826
rect 3570 -2860 3604 -2826
rect 3638 -2860 3672 -2826
rect 3706 -2860 3850 -2826
rect 3884 -2860 3918 -2826
rect 3952 -2860 3986 -2826
rect 4020 -2860 4054 -2826
rect 4088 -2860 4288 -2826
rect 4322 -2860 4356 -2826
rect 4390 -2860 4424 -2826
rect 4458 -2860 4492 -2826
rect 4526 -2860 4670 -2826
rect 4704 -2860 4738 -2826
rect 4772 -2860 4806 -2826
rect 4840 -2860 4874 -2826
rect 4908 -2860 5108 -2826
rect 5142 -2860 5176 -2826
rect 5210 -2860 5244 -2826
rect 5278 -2860 5312 -2826
rect 5346 -2860 5490 -2826
rect 5524 -2860 5558 -2826
rect 5592 -2860 5626 -2826
rect 5660 -2860 5694 -2826
rect 5728 -2860 5928 -2826
rect 5962 -2860 5996 -2826
rect 6030 -2860 6064 -2826
rect 6098 -2860 6132 -2826
rect 6166 -2860 6310 -2826
rect 6344 -2860 6378 -2826
rect 6412 -2860 6446 -2826
rect 6480 -2860 6514 -2826
rect 6548 -2860 6748 -2826
rect 6782 -2860 6816 -2826
rect 6850 -2860 6884 -2826
rect 6918 -2860 6952 -2826
rect 6986 -2860 7030 -2826
rect -1110 -3004 7030 -2860
rect -1110 -3038 -1070 -3004
rect -1036 -3038 -1002 -3004
rect -968 -3038 -934 -3004
rect -900 -3038 -866 -3004
rect -832 -3038 -632 -3004
rect -598 -3038 -564 -3004
rect -530 -3038 -496 -3004
rect -462 -3038 -428 -3004
rect -394 -3038 -250 -3004
rect -216 -3038 -182 -3004
rect -148 -3038 -114 -3004
rect -80 -3038 -46 -3004
rect -12 -3038 188 -3004
rect 222 -3038 256 -3004
rect 290 -3038 324 -3004
rect 358 -3038 392 -3004
rect 426 -3038 570 -3004
rect 604 -3038 638 -3004
rect 672 -3038 706 -3004
rect 740 -3038 774 -3004
rect 808 -3038 1008 -3004
rect 1042 -3038 1076 -3004
rect 1110 -3038 1144 -3004
rect 1178 -3038 1212 -3004
rect 1246 -3038 1390 -3004
rect 1424 -3038 1458 -3004
rect 1492 -3038 1526 -3004
rect 1560 -3038 1594 -3004
rect 1628 -3038 1828 -3004
rect 1862 -3038 1896 -3004
rect 1930 -3038 1964 -3004
rect 1998 -3038 2032 -3004
rect 2066 -3038 2210 -3004
rect 2244 -3038 2278 -3004
rect 2312 -3038 2346 -3004
rect 2380 -3038 2414 -3004
rect 2448 -3038 2648 -3004
rect 2682 -3038 2716 -3004
rect 2750 -3038 2784 -3004
rect 2818 -3038 2852 -3004
rect 2886 -3038 3030 -3004
rect 3064 -3038 3098 -3004
rect 3132 -3038 3166 -3004
rect 3200 -3038 3234 -3004
rect 3268 -3038 3468 -3004
rect 3502 -3038 3536 -3004
rect 3570 -3038 3604 -3004
rect 3638 -3038 3672 -3004
rect 3706 -3038 3850 -3004
rect 3884 -3038 3918 -3004
rect 3952 -3038 3986 -3004
rect 4020 -3038 4054 -3004
rect 4088 -3038 4288 -3004
rect 4322 -3038 4356 -3004
rect 4390 -3038 4424 -3004
rect 4458 -3038 4492 -3004
rect 4526 -3038 4670 -3004
rect 4704 -3038 4738 -3004
rect 4772 -3038 4806 -3004
rect 4840 -3038 4874 -3004
rect 4908 -3038 5108 -3004
rect 5142 -3038 5176 -3004
rect 5210 -3038 5244 -3004
rect 5278 -3038 5312 -3004
rect 5346 -3038 5490 -3004
rect 5524 -3038 5558 -3004
rect 5592 -3038 5626 -3004
rect 5660 -3038 5694 -3004
rect 5728 -3038 5928 -3004
rect 5962 -3038 5996 -3004
rect 6030 -3038 6064 -3004
rect 6098 -3038 6132 -3004
rect 6166 -3038 6310 -3004
rect 6344 -3038 6378 -3004
rect 6412 -3038 6446 -3004
rect 6480 -3038 6514 -3004
rect 6548 -3038 6748 -3004
rect 6782 -3038 6816 -3004
rect 6850 -3038 6884 -3004
rect 6918 -3038 6952 -3004
rect 6986 -3038 7030 -3004
rect -1110 -3072 7030 -3038
rect -1110 -3106 -1070 -3072
rect -1036 -3106 -428 -3072
rect -394 -3106 -250 -3072
rect -216 -3106 392 -3072
rect 426 -3106 570 -3072
rect 604 -3106 1212 -3072
rect 1246 -3106 1390 -3072
rect 1424 -3106 2032 -3072
rect 2066 -3106 2210 -3072
rect 2244 -3106 2852 -3072
rect 2886 -3106 3030 -3072
rect 3064 -3106 3672 -3072
rect 3706 -3106 3850 -3072
rect 3884 -3106 4492 -3072
rect 4526 -3106 4670 -3072
rect 4704 -3106 5312 -3072
rect 5346 -3106 5490 -3072
rect 5524 -3106 6132 -3072
rect 6166 -3106 6310 -3072
rect 6344 -3106 6952 -3072
rect 6986 -3106 7030 -3072
rect -1110 -3140 7030 -3106
rect -1110 -3174 -1070 -3140
rect -1036 -3157 -428 -3140
rect -1036 -3174 -917 -3157
rect -1110 -3191 -917 -3174
rect -883 -3191 -849 -3157
rect -815 -3191 -649 -3157
rect -615 -3191 -581 -3157
rect -547 -3174 -428 -3157
rect -394 -3174 -250 -3140
rect -216 -3157 392 -3140
rect -216 -3174 -97 -3157
rect -547 -3191 -97 -3174
rect -63 -3191 -29 -3157
rect 5 -3191 171 -3157
rect 205 -3191 239 -3157
rect 273 -3174 392 -3157
rect 426 -3174 570 -3140
rect 604 -3157 1212 -3140
rect 604 -3174 723 -3157
rect 273 -3191 723 -3174
rect 757 -3191 791 -3157
rect 825 -3191 991 -3157
rect 1025 -3191 1059 -3157
rect 1093 -3174 1212 -3157
rect 1246 -3174 1390 -3140
rect 1424 -3157 2032 -3140
rect 1424 -3174 1543 -3157
rect 1093 -3191 1543 -3174
rect 1577 -3191 1611 -3157
rect 1645 -3191 1811 -3157
rect 1845 -3191 1879 -3157
rect 1913 -3174 2032 -3157
rect 2066 -3174 2210 -3140
rect 2244 -3157 2852 -3140
rect 2244 -3174 2363 -3157
rect 1913 -3191 2363 -3174
rect 2397 -3191 2431 -3157
rect 2465 -3191 2631 -3157
rect 2665 -3191 2699 -3157
rect 2733 -3174 2852 -3157
rect 2886 -3174 3030 -3140
rect 3064 -3157 3672 -3140
rect 3064 -3174 3183 -3157
rect 2733 -3191 3183 -3174
rect 3217 -3191 3251 -3157
rect 3285 -3191 3451 -3157
rect 3485 -3191 3519 -3157
rect 3553 -3174 3672 -3157
rect 3706 -3174 3850 -3140
rect 3884 -3157 4492 -3140
rect 3884 -3174 4003 -3157
rect 3553 -3191 4003 -3174
rect 4037 -3191 4071 -3157
rect 4105 -3191 4271 -3157
rect 4305 -3191 4339 -3157
rect 4373 -3174 4492 -3157
rect 4526 -3174 4670 -3140
rect 4704 -3157 5312 -3140
rect 4704 -3174 4823 -3157
rect 4373 -3191 4823 -3174
rect 4857 -3191 4891 -3157
rect 4925 -3191 5091 -3157
rect 5125 -3191 5159 -3157
rect 5193 -3174 5312 -3157
rect 5346 -3174 5490 -3140
rect 5524 -3157 6132 -3140
rect 5524 -3174 5643 -3157
rect 5193 -3191 5643 -3174
rect 5677 -3191 5711 -3157
rect 5745 -3191 5911 -3157
rect 5945 -3191 5979 -3157
rect 6013 -3174 6132 -3157
rect 6166 -3174 6310 -3140
rect 6344 -3157 6952 -3140
rect 6344 -3174 6463 -3157
rect 6013 -3191 6463 -3174
rect 6497 -3191 6531 -3157
rect 6565 -3191 6731 -3157
rect 6765 -3191 6799 -3157
rect 6833 -3174 6952 -3157
rect 6986 -3174 7030 -3140
rect 6833 -3191 7030 -3174
rect 15940 -3180 16190 -2740
rect -1110 -3208 7030 -3191
rect -1110 -3210 -1070 -3208
rect -1104 -3242 -1070 -3210
rect -1036 -3210 -428 -3208
rect -1036 -3242 -1003 -3210
rect -1104 -3442 -1003 -3242
rect -1104 -3470 -1070 -3442
rect -1110 -3476 -1070 -3470
rect -1036 -3470 -1003 -3442
rect -941 -3225 -869 -3210
rect -941 -3259 -917 -3225
rect -883 -3259 -869 -3225
rect -941 -3425 -869 -3259
rect -595 -3225 -523 -3210
rect -595 -3259 -581 -3225
rect -547 -3259 -523 -3225
rect -811 -3277 -653 -3263
rect -811 -3311 -797 -3277
rect -763 -3291 -701 -3277
rect -667 -3311 -653 -3277
rect -811 -3373 -783 -3311
rect -681 -3373 -653 -3311
rect -811 -3407 -797 -3373
rect -763 -3407 -701 -3393
rect -667 -3407 -653 -3373
rect -811 -3421 -653 -3407
rect -941 -3459 -917 -3425
rect -883 -3459 -869 -3425
rect -941 -3470 -869 -3459
rect -595 -3425 -523 -3259
rect -595 -3459 -581 -3425
rect -547 -3459 -523 -3425
rect -595 -3470 -523 -3459
rect -461 -3242 -428 -3210
rect -394 -3210 -250 -3208
rect -394 -3242 -360 -3210
rect -461 -3442 -360 -3242
rect -461 -3470 -428 -3442
rect -1036 -3476 -428 -3470
rect -394 -3470 -360 -3442
rect -284 -3242 -250 -3210
rect -216 -3210 392 -3208
rect -216 -3242 -183 -3210
rect -284 -3442 -183 -3242
rect -284 -3470 -250 -3442
rect -394 -3476 -250 -3470
rect -216 -3470 -183 -3442
rect -121 -3225 -49 -3210
rect -121 -3259 -97 -3225
rect -63 -3259 -49 -3225
rect -121 -3425 -49 -3259
rect 225 -3225 297 -3210
rect 225 -3259 239 -3225
rect 273 -3259 297 -3225
rect 9 -3277 167 -3263
rect 9 -3311 23 -3277
rect 57 -3291 119 -3277
rect 153 -3311 167 -3277
rect 9 -3373 37 -3311
rect 139 -3373 167 -3311
rect 9 -3407 23 -3373
rect 57 -3407 119 -3393
rect 153 -3407 167 -3373
rect 9 -3421 167 -3407
rect -121 -3459 -97 -3425
rect -63 -3459 -49 -3425
rect -121 -3470 -49 -3459
rect 225 -3425 297 -3259
rect 225 -3459 239 -3425
rect 273 -3459 297 -3425
rect 225 -3470 297 -3459
rect 359 -3242 392 -3210
rect 426 -3210 570 -3208
rect 426 -3242 460 -3210
rect 359 -3442 460 -3242
rect 359 -3470 392 -3442
rect -216 -3476 392 -3470
rect 426 -3470 460 -3442
rect 536 -3242 570 -3210
rect 604 -3210 1212 -3208
rect 604 -3242 637 -3210
rect 536 -3442 637 -3242
rect 536 -3470 570 -3442
rect 426 -3476 570 -3470
rect 604 -3470 637 -3442
rect 699 -3225 771 -3210
rect 699 -3259 723 -3225
rect 757 -3259 771 -3225
rect 699 -3425 771 -3259
rect 1045 -3225 1117 -3210
rect 1045 -3259 1059 -3225
rect 1093 -3259 1117 -3225
rect 829 -3277 987 -3263
rect 829 -3311 843 -3277
rect 877 -3291 939 -3277
rect 973 -3311 987 -3277
rect 829 -3373 857 -3311
rect 959 -3373 987 -3311
rect 829 -3407 843 -3373
rect 877 -3407 939 -3393
rect 973 -3407 987 -3373
rect 829 -3421 987 -3407
rect 699 -3459 723 -3425
rect 757 -3459 771 -3425
rect 699 -3470 771 -3459
rect 1045 -3425 1117 -3259
rect 1045 -3459 1059 -3425
rect 1093 -3459 1117 -3425
rect 1045 -3470 1117 -3459
rect 1179 -3242 1212 -3210
rect 1246 -3210 1390 -3208
rect 1246 -3242 1280 -3210
rect 1179 -3442 1280 -3242
rect 1179 -3470 1212 -3442
rect 604 -3476 1212 -3470
rect 1246 -3470 1280 -3442
rect 1356 -3242 1390 -3210
rect 1424 -3210 2032 -3208
rect 1424 -3242 1457 -3210
rect 1356 -3442 1457 -3242
rect 1356 -3470 1390 -3442
rect 1246 -3476 1390 -3470
rect 1424 -3470 1457 -3442
rect 1519 -3225 1591 -3210
rect 1519 -3259 1543 -3225
rect 1577 -3259 1591 -3225
rect 1519 -3425 1591 -3259
rect 1865 -3225 1937 -3210
rect 1865 -3259 1879 -3225
rect 1913 -3259 1937 -3225
rect 1649 -3277 1807 -3263
rect 1649 -3311 1663 -3277
rect 1697 -3291 1759 -3277
rect 1793 -3311 1807 -3277
rect 1649 -3373 1677 -3311
rect 1779 -3373 1807 -3311
rect 1649 -3407 1663 -3373
rect 1697 -3407 1759 -3393
rect 1793 -3407 1807 -3373
rect 1649 -3421 1807 -3407
rect 1519 -3459 1543 -3425
rect 1577 -3459 1591 -3425
rect 1519 -3470 1591 -3459
rect 1865 -3425 1937 -3259
rect 1865 -3459 1879 -3425
rect 1913 -3459 1937 -3425
rect 1865 -3470 1937 -3459
rect 1999 -3242 2032 -3210
rect 2066 -3210 2210 -3208
rect 2066 -3242 2100 -3210
rect 1999 -3442 2100 -3242
rect 1999 -3470 2032 -3442
rect 1424 -3476 2032 -3470
rect 2066 -3470 2100 -3442
rect 2176 -3242 2210 -3210
rect 2244 -3210 2852 -3208
rect 2244 -3242 2277 -3210
rect 2176 -3442 2277 -3242
rect 2176 -3470 2210 -3442
rect 2066 -3476 2210 -3470
rect 2244 -3470 2277 -3442
rect 2339 -3225 2411 -3210
rect 2339 -3259 2363 -3225
rect 2397 -3259 2411 -3225
rect 2339 -3425 2411 -3259
rect 2685 -3225 2757 -3210
rect 2685 -3259 2699 -3225
rect 2733 -3259 2757 -3225
rect 2469 -3277 2627 -3263
rect 2469 -3311 2483 -3277
rect 2517 -3291 2579 -3277
rect 2613 -3311 2627 -3277
rect 2469 -3373 2497 -3311
rect 2599 -3373 2627 -3311
rect 2469 -3407 2483 -3373
rect 2517 -3407 2579 -3393
rect 2613 -3407 2627 -3373
rect 2469 -3421 2627 -3407
rect 2339 -3459 2363 -3425
rect 2397 -3459 2411 -3425
rect 2339 -3470 2411 -3459
rect 2685 -3425 2757 -3259
rect 2685 -3459 2699 -3425
rect 2733 -3459 2757 -3425
rect 2685 -3470 2757 -3459
rect 2819 -3242 2852 -3210
rect 2886 -3210 3030 -3208
rect 2886 -3242 2920 -3210
rect 2819 -3442 2920 -3242
rect 2819 -3470 2852 -3442
rect 2244 -3476 2852 -3470
rect 2886 -3470 2920 -3442
rect 2996 -3242 3030 -3210
rect 3064 -3210 3672 -3208
rect 3064 -3242 3097 -3210
rect 2996 -3442 3097 -3242
rect 2996 -3470 3030 -3442
rect 2886 -3476 3030 -3470
rect 3064 -3470 3097 -3442
rect 3159 -3225 3231 -3210
rect 3159 -3259 3183 -3225
rect 3217 -3259 3231 -3225
rect 3159 -3425 3231 -3259
rect 3505 -3225 3577 -3210
rect 3505 -3259 3519 -3225
rect 3553 -3259 3577 -3225
rect 3289 -3277 3447 -3263
rect 3289 -3311 3303 -3277
rect 3337 -3291 3399 -3277
rect 3433 -3311 3447 -3277
rect 3289 -3373 3317 -3311
rect 3419 -3373 3447 -3311
rect 3289 -3407 3303 -3373
rect 3337 -3407 3399 -3393
rect 3433 -3407 3447 -3373
rect 3289 -3421 3447 -3407
rect 3159 -3459 3183 -3425
rect 3217 -3459 3231 -3425
rect 3159 -3470 3231 -3459
rect 3505 -3425 3577 -3259
rect 3505 -3459 3519 -3425
rect 3553 -3459 3577 -3425
rect 3505 -3470 3577 -3459
rect 3639 -3242 3672 -3210
rect 3706 -3210 3850 -3208
rect 3706 -3242 3740 -3210
rect 3639 -3442 3740 -3242
rect 3639 -3470 3672 -3442
rect 3064 -3476 3672 -3470
rect 3706 -3470 3740 -3442
rect 3816 -3242 3850 -3210
rect 3884 -3210 4492 -3208
rect 3884 -3242 3917 -3210
rect 3816 -3442 3917 -3242
rect 3816 -3470 3850 -3442
rect 3706 -3476 3850 -3470
rect 3884 -3470 3917 -3442
rect 3979 -3225 4051 -3210
rect 3979 -3259 4003 -3225
rect 4037 -3259 4051 -3225
rect 3979 -3425 4051 -3259
rect 4325 -3225 4397 -3210
rect 4325 -3259 4339 -3225
rect 4373 -3259 4397 -3225
rect 4109 -3277 4267 -3263
rect 4109 -3311 4123 -3277
rect 4157 -3291 4219 -3277
rect 4253 -3311 4267 -3277
rect 4109 -3373 4137 -3311
rect 4239 -3373 4267 -3311
rect 4109 -3407 4123 -3373
rect 4157 -3407 4219 -3393
rect 4253 -3407 4267 -3373
rect 4109 -3421 4267 -3407
rect 3979 -3459 4003 -3425
rect 4037 -3459 4051 -3425
rect 3979 -3470 4051 -3459
rect 4325 -3425 4397 -3259
rect 4325 -3459 4339 -3425
rect 4373 -3459 4397 -3425
rect 4325 -3470 4397 -3459
rect 4459 -3242 4492 -3210
rect 4526 -3210 4670 -3208
rect 4526 -3242 4560 -3210
rect 4459 -3442 4560 -3242
rect 4459 -3470 4492 -3442
rect 3884 -3476 4492 -3470
rect 4526 -3470 4560 -3442
rect 4636 -3242 4670 -3210
rect 4704 -3210 5312 -3208
rect 4704 -3242 4737 -3210
rect 4636 -3442 4737 -3242
rect 4636 -3470 4670 -3442
rect 4526 -3476 4670 -3470
rect 4704 -3470 4737 -3442
rect 4799 -3225 4871 -3210
rect 4799 -3259 4823 -3225
rect 4857 -3259 4871 -3225
rect 4799 -3425 4871 -3259
rect 5145 -3225 5217 -3210
rect 5145 -3259 5159 -3225
rect 5193 -3259 5217 -3225
rect 4929 -3277 5087 -3263
rect 4929 -3311 4943 -3277
rect 4977 -3291 5039 -3277
rect 5073 -3311 5087 -3277
rect 4929 -3373 4957 -3311
rect 5059 -3373 5087 -3311
rect 4929 -3407 4943 -3373
rect 4977 -3407 5039 -3393
rect 5073 -3407 5087 -3373
rect 4929 -3421 5087 -3407
rect 4799 -3459 4823 -3425
rect 4857 -3459 4871 -3425
rect 4799 -3470 4871 -3459
rect 5145 -3425 5217 -3259
rect 5145 -3459 5159 -3425
rect 5193 -3459 5217 -3425
rect 5145 -3470 5217 -3459
rect 5279 -3242 5312 -3210
rect 5346 -3210 5490 -3208
rect 5346 -3242 5380 -3210
rect 5279 -3442 5380 -3242
rect 5279 -3470 5312 -3442
rect 4704 -3476 5312 -3470
rect 5346 -3470 5380 -3442
rect 5456 -3242 5490 -3210
rect 5524 -3210 6132 -3208
rect 5524 -3242 5557 -3210
rect 5456 -3442 5557 -3242
rect 5456 -3470 5490 -3442
rect 5346 -3476 5490 -3470
rect 5524 -3470 5557 -3442
rect 5619 -3225 5691 -3210
rect 5619 -3259 5643 -3225
rect 5677 -3259 5691 -3225
rect 5619 -3425 5691 -3259
rect 5965 -3225 6037 -3210
rect 5965 -3259 5979 -3225
rect 6013 -3259 6037 -3225
rect 5749 -3277 5907 -3263
rect 5749 -3311 5763 -3277
rect 5797 -3291 5859 -3277
rect 5893 -3311 5907 -3277
rect 5749 -3373 5777 -3311
rect 5879 -3373 5907 -3311
rect 5749 -3407 5763 -3373
rect 5797 -3407 5859 -3393
rect 5893 -3407 5907 -3373
rect 5749 -3421 5907 -3407
rect 5619 -3459 5643 -3425
rect 5677 -3459 5691 -3425
rect 5619 -3470 5691 -3459
rect 5965 -3425 6037 -3259
rect 5965 -3459 5979 -3425
rect 6013 -3459 6037 -3425
rect 5965 -3470 6037 -3459
rect 6099 -3242 6132 -3210
rect 6166 -3210 6310 -3208
rect 6166 -3242 6200 -3210
rect 6099 -3442 6200 -3242
rect 6099 -3470 6132 -3442
rect 5524 -3476 6132 -3470
rect 6166 -3470 6200 -3442
rect 6276 -3242 6310 -3210
rect 6344 -3210 6952 -3208
rect 6344 -3242 6377 -3210
rect 6276 -3442 6377 -3242
rect 6276 -3470 6310 -3442
rect 6166 -3476 6310 -3470
rect 6344 -3470 6377 -3442
rect 6439 -3225 6511 -3210
rect 6439 -3259 6463 -3225
rect 6497 -3259 6511 -3225
rect 6439 -3425 6511 -3259
rect 6785 -3225 6857 -3210
rect 6785 -3259 6799 -3225
rect 6833 -3259 6857 -3225
rect 6569 -3277 6727 -3263
rect 6569 -3311 6583 -3277
rect 6617 -3291 6679 -3277
rect 6713 -3311 6727 -3277
rect 6569 -3373 6597 -3311
rect 6699 -3373 6727 -3311
rect 6569 -3407 6583 -3373
rect 6617 -3407 6679 -3393
rect 6713 -3407 6727 -3373
rect 6569 -3421 6727 -3407
rect 6439 -3459 6463 -3425
rect 6497 -3459 6511 -3425
rect 6439 -3470 6511 -3459
rect 6785 -3425 6857 -3259
rect 6785 -3459 6799 -3425
rect 6833 -3459 6857 -3425
rect 6785 -3470 6857 -3459
rect 6919 -3242 6952 -3210
rect 6986 -3210 7030 -3208
rect 6986 -3242 7020 -3210
rect 16410 -3240 16500 -1340
rect 16720 -3180 16970 -2740
rect 6919 -3442 7020 -3242
rect 6919 -3470 6952 -3442
rect 6344 -3476 6952 -3470
rect 6986 -3470 7020 -3442
rect 15760 -3320 16500 -3240
rect 6986 -3476 7030 -3470
rect -1110 -3493 7030 -3476
rect -1110 -3510 -917 -3493
rect -1110 -3544 -1070 -3510
rect -1036 -3527 -917 -3510
rect -883 -3527 -849 -3493
rect -815 -3527 -649 -3493
rect -615 -3527 -581 -3493
rect -547 -3510 -97 -3493
rect -547 -3527 -428 -3510
rect -1036 -3544 -428 -3527
rect -394 -3544 -250 -3510
rect -216 -3527 -97 -3510
rect -63 -3527 -29 -3493
rect 5 -3527 171 -3493
rect 205 -3527 239 -3493
rect 273 -3510 723 -3493
rect 273 -3527 392 -3510
rect -216 -3544 392 -3527
rect 426 -3544 570 -3510
rect 604 -3527 723 -3510
rect 757 -3527 791 -3493
rect 825 -3527 991 -3493
rect 1025 -3527 1059 -3493
rect 1093 -3510 1543 -3493
rect 1093 -3527 1212 -3510
rect 604 -3544 1212 -3527
rect 1246 -3544 1390 -3510
rect 1424 -3527 1543 -3510
rect 1577 -3527 1611 -3493
rect 1645 -3527 1811 -3493
rect 1845 -3527 1879 -3493
rect 1913 -3510 2363 -3493
rect 1913 -3527 2032 -3510
rect 1424 -3544 2032 -3527
rect 2066 -3544 2210 -3510
rect 2244 -3527 2363 -3510
rect 2397 -3527 2431 -3493
rect 2465 -3527 2631 -3493
rect 2665 -3527 2699 -3493
rect 2733 -3510 3183 -3493
rect 2733 -3527 2852 -3510
rect 2244 -3544 2852 -3527
rect 2886 -3544 3030 -3510
rect 3064 -3527 3183 -3510
rect 3217 -3527 3251 -3493
rect 3285 -3527 3451 -3493
rect 3485 -3527 3519 -3493
rect 3553 -3510 4003 -3493
rect 3553 -3527 3672 -3510
rect 3064 -3544 3672 -3527
rect 3706 -3544 3850 -3510
rect 3884 -3527 4003 -3510
rect 4037 -3527 4071 -3493
rect 4105 -3527 4271 -3493
rect 4305 -3527 4339 -3493
rect 4373 -3510 4823 -3493
rect 4373 -3527 4492 -3510
rect 3884 -3544 4492 -3527
rect 4526 -3544 4670 -3510
rect 4704 -3527 4823 -3510
rect 4857 -3527 4891 -3493
rect 4925 -3527 5091 -3493
rect 5125 -3527 5159 -3493
rect 5193 -3510 5643 -3493
rect 5193 -3527 5312 -3510
rect 4704 -3544 5312 -3527
rect 5346 -3544 5490 -3510
rect 5524 -3527 5643 -3510
rect 5677 -3527 5711 -3493
rect 5745 -3527 5911 -3493
rect 5945 -3527 5979 -3493
rect 6013 -3510 6463 -3493
rect 6013 -3527 6132 -3510
rect 5524 -3544 6132 -3527
rect 6166 -3544 6310 -3510
rect 6344 -3527 6463 -3510
rect 6497 -3527 6531 -3493
rect 6565 -3527 6731 -3493
rect 6765 -3527 6799 -3493
rect 6833 -3510 7030 -3493
rect 6833 -3527 6952 -3510
rect 6344 -3544 6952 -3527
rect 6986 -3544 7030 -3510
rect -1110 -3578 7030 -3544
rect -1110 -3612 -1070 -3578
rect -1036 -3612 -428 -3578
rect -394 -3612 -250 -3578
rect -216 -3612 392 -3578
rect 426 -3612 570 -3578
rect 604 -3612 1212 -3578
rect 1246 -3612 1390 -3578
rect 1424 -3612 2032 -3578
rect 2066 -3612 2210 -3578
rect 2244 -3612 2852 -3578
rect 2886 -3612 3030 -3578
rect 3064 -3612 3672 -3578
rect 3706 -3612 3850 -3578
rect 3884 -3612 4492 -3578
rect 4526 -3612 4670 -3578
rect 4704 -3612 5312 -3578
rect 5346 -3612 5490 -3578
rect 5524 -3612 6132 -3578
rect 6166 -3612 6310 -3578
rect 6344 -3612 6952 -3578
rect 6986 -3612 7030 -3578
rect -1110 -3646 7030 -3612
rect -1110 -3680 -1070 -3646
rect -1036 -3680 -1002 -3646
rect -968 -3680 -934 -3646
rect -900 -3680 -866 -3646
rect -832 -3680 -632 -3646
rect -598 -3680 -564 -3646
rect -530 -3680 -496 -3646
rect -462 -3680 -428 -3646
rect -394 -3680 -250 -3646
rect -216 -3680 -182 -3646
rect -148 -3680 -114 -3646
rect -80 -3680 -46 -3646
rect -12 -3680 188 -3646
rect 222 -3680 256 -3646
rect 290 -3680 324 -3646
rect 358 -3680 392 -3646
rect 426 -3680 570 -3646
rect 604 -3680 638 -3646
rect 672 -3680 706 -3646
rect 740 -3680 774 -3646
rect 808 -3680 1008 -3646
rect 1042 -3680 1076 -3646
rect 1110 -3680 1144 -3646
rect 1178 -3680 1212 -3646
rect 1246 -3680 1390 -3646
rect 1424 -3680 1458 -3646
rect 1492 -3680 1526 -3646
rect 1560 -3680 1594 -3646
rect 1628 -3680 1828 -3646
rect 1862 -3680 1896 -3646
rect 1930 -3680 1964 -3646
rect 1998 -3680 2032 -3646
rect 2066 -3680 2210 -3646
rect 2244 -3680 2278 -3646
rect 2312 -3680 2346 -3646
rect 2380 -3680 2414 -3646
rect 2448 -3680 2648 -3646
rect 2682 -3680 2716 -3646
rect 2750 -3680 2784 -3646
rect 2818 -3680 2852 -3646
rect 2886 -3680 3030 -3646
rect 3064 -3680 3098 -3646
rect 3132 -3680 3166 -3646
rect 3200 -3680 3234 -3646
rect 3268 -3680 3468 -3646
rect 3502 -3680 3536 -3646
rect 3570 -3680 3604 -3646
rect 3638 -3680 3672 -3646
rect 3706 -3680 3850 -3646
rect 3884 -3680 3918 -3646
rect 3952 -3680 3986 -3646
rect 4020 -3680 4054 -3646
rect 4088 -3680 4288 -3646
rect 4322 -3680 4356 -3646
rect 4390 -3680 4424 -3646
rect 4458 -3680 4492 -3646
rect 4526 -3680 4670 -3646
rect 4704 -3680 4738 -3646
rect 4772 -3680 4806 -3646
rect 4840 -3680 4874 -3646
rect 4908 -3680 5108 -3646
rect 5142 -3680 5176 -3646
rect 5210 -3680 5244 -3646
rect 5278 -3680 5312 -3646
rect 5346 -3680 5490 -3646
rect 5524 -3680 5558 -3646
rect 5592 -3680 5626 -3646
rect 5660 -3680 5694 -3646
rect 5728 -3680 5928 -3646
rect 5962 -3680 5996 -3646
rect 6030 -3680 6064 -3646
rect 6098 -3680 6132 -3646
rect 6166 -3680 6310 -3646
rect 6344 -3680 6378 -3646
rect 6412 -3680 6446 -3646
rect 6480 -3680 6514 -3646
rect 6548 -3680 6748 -3646
rect 6782 -3680 6816 -3646
rect 6850 -3680 6884 -3646
rect 6918 -3680 6952 -3646
rect 6986 -3680 7030 -3646
rect -1110 -3824 7030 -3680
rect -1110 -3858 -1070 -3824
rect -1036 -3858 -1002 -3824
rect -968 -3858 -934 -3824
rect -900 -3858 -866 -3824
rect -832 -3858 -632 -3824
rect -598 -3858 -564 -3824
rect -530 -3858 -496 -3824
rect -462 -3858 -428 -3824
rect -394 -3858 -250 -3824
rect -216 -3858 -182 -3824
rect -148 -3858 -114 -3824
rect -80 -3858 -46 -3824
rect -12 -3858 188 -3824
rect 222 -3858 256 -3824
rect 290 -3858 324 -3824
rect 358 -3858 392 -3824
rect 426 -3858 570 -3824
rect 604 -3858 638 -3824
rect 672 -3858 706 -3824
rect 740 -3858 774 -3824
rect 808 -3858 1008 -3824
rect 1042 -3858 1076 -3824
rect 1110 -3858 1144 -3824
rect 1178 -3858 1212 -3824
rect 1246 -3858 1390 -3824
rect 1424 -3858 1458 -3824
rect 1492 -3858 1526 -3824
rect 1560 -3858 1594 -3824
rect 1628 -3858 1828 -3824
rect 1862 -3858 1896 -3824
rect 1930 -3858 1964 -3824
rect 1998 -3858 2032 -3824
rect 2066 -3858 2210 -3824
rect 2244 -3858 2278 -3824
rect 2312 -3858 2346 -3824
rect 2380 -3858 2414 -3824
rect 2448 -3858 2648 -3824
rect 2682 -3858 2716 -3824
rect 2750 -3858 2784 -3824
rect 2818 -3858 2852 -3824
rect 2886 -3858 3030 -3824
rect 3064 -3858 3098 -3824
rect 3132 -3858 3166 -3824
rect 3200 -3858 3234 -3824
rect 3268 -3858 3468 -3824
rect 3502 -3858 3536 -3824
rect 3570 -3858 3604 -3824
rect 3638 -3858 3672 -3824
rect 3706 -3858 3850 -3824
rect 3884 -3858 3918 -3824
rect 3952 -3858 3986 -3824
rect 4020 -3858 4054 -3824
rect 4088 -3858 4288 -3824
rect 4322 -3858 4356 -3824
rect 4390 -3858 4424 -3824
rect 4458 -3858 4492 -3824
rect 4526 -3858 4670 -3824
rect 4704 -3858 4738 -3824
rect 4772 -3858 4806 -3824
rect 4840 -3858 4874 -3824
rect 4908 -3858 5108 -3824
rect 5142 -3858 5176 -3824
rect 5210 -3858 5244 -3824
rect 5278 -3858 5312 -3824
rect 5346 -3858 5490 -3824
rect 5524 -3858 5558 -3824
rect 5592 -3858 5626 -3824
rect 5660 -3858 5694 -3824
rect 5728 -3858 5928 -3824
rect 5962 -3858 5996 -3824
rect 6030 -3858 6064 -3824
rect 6098 -3858 6132 -3824
rect 6166 -3858 6310 -3824
rect 6344 -3858 6378 -3824
rect 6412 -3858 6446 -3824
rect 6480 -3858 6514 -3824
rect 6548 -3858 6748 -3824
rect 6782 -3858 6816 -3824
rect 6850 -3858 6884 -3824
rect 6918 -3858 6952 -3824
rect 6986 -3858 7030 -3824
rect -1110 -3892 7030 -3858
rect -1110 -3926 -1070 -3892
rect -1036 -3926 -428 -3892
rect -394 -3926 -250 -3892
rect -216 -3926 392 -3892
rect 426 -3926 570 -3892
rect 604 -3926 1212 -3892
rect 1246 -3926 1390 -3892
rect 1424 -3926 2032 -3892
rect 2066 -3926 2210 -3892
rect 2244 -3926 2852 -3892
rect 2886 -3926 3030 -3892
rect 3064 -3926 3672 -3892
rect 3706 -3926 3850 -3892
rect 3884 -3926 4492 -3892
rect 4526 -3926 4670 -3892
rect 4704 -3926 5312 -3892
rect 5346 -3926 5490 -3892
rect 5524 -3926 6132 -3892
rect 6166 -3926 6310 -3892
rect 6344 -3926 6952 -3892
rect 6986 -3926 7030 -3892
rect -1110 -3960 7030 -3926
rect -1110 -3994 -1070 -3960
rect -1036 -3977 -428 -3960
rect -1036 -3994 -917 -3977
rect -1110 -4011 -917 -3994
rect -883 -4011 -849 -3977
rect -815 -4011 -649 -3977
rect -615 -4011 -581 -3977
rect -547 -3994 -428 -3977
rect -394 -3994 -250 -3960
rect -216 -3977 392 -3960
rect -216 -3994 -97 -3977
rect -547 -4011 -97 -3994
rect -63 -4011 -29 -3977
rect 5 -4011 171 -3977
rect 205 -4011 239 -3977
rect 273 -3994 392 -3977
rect 426 -3994 570 -3960
rect 604 -3977 1212 -3960
rect 604 -3994 723 -3977
rect 273 -4011 723 -3994
rect 757 -4011 791 -3977
rect 825 -4011 991 -3977
rect 1025 -4011 1059 -3977
rect 1093 -3994 1212 -3977
rect 1246 -3994 1390 -3960
rect 1424 -3977 2032 -3960
rect 1424 -3994 1543 -3977
rect 1093 -4011 1543 -3994
rect 1577 -4011 1611 -3977
rect 1645 -4011 1811 -3977
rect 1845 -4011 1879 -3977
rect 1913 -3994 2032 -3977
rect 2066 -3994 2210 -3960
rect 2244 -3977 2852 -3960
rect 2244 -3994 2363 -3977
rect 1913 -4011 2363 -3994
rect 2397 -4011 2431 -3977
rect 2465 -4011 2631 -3977
rect 2665 -4011 2699 -3977
rect 2733 -3994 2852 -3977
rect 2886 -3994 3030 -3960
rect 3064 -3977 3672 -3960
rect 3064 -3994 3183 -3977
rect 2733 -4011 3183 -3994
rect 3217 -4011 3251 -3977
rect 3285 -4011 3451 -3977
rect 3485 -4011 3519 -3977
rect 3553 -3994 3672 -3977
rect 3706 -3994 3850 -3960
rect 3884 -3977 4492 -3960
rect 3884 -3994 4003 -3977
rect 3553 -4011 4003 -3994
rect 4037 -4011 4071 -3977
rect 4105 -4011 4271 -3977
rect 4305 -4011 4339 -3977
rect 4373 -3994 4492 -3977
rect 4526 -3994 4670 -3960
rect 4704 -3977 5312 -3960
rect 4704 -3994 4823 -3977
rect 4373 -4011 4823 -3994
rect 4857 -4011 4891 -3977
rect 4925 -4011 5091 -3977
rect 5125 -4011 5159 -3977
rect 5193 -3994 5312 -3977
rect 5346 -3994 5490 -3960
rect 5524 -3977 6132 -3960
rect 5524 -3994 5643 -3977
rect 5193 -4011 5643 -3994
rect 5677 -4011 5711 -3977
rect 5745 -4011 5911 -3977
rect 5945 -4011 5979 -3977
rect 6013 -3994 6132 -3977
rect 6166 -3994 6310 -3960
rect 6344 -3977 6952 -3960
rect 6344 -3994 6463 -3977
rect 6013 -4011 6463 -3994
rect 6497 -4011 6531 -3977
rect 6565 -4011 6731 -3977
rect 6765 -4011 6799 -3977
rect 6833 -3994 6952 -3977
rect 6986 -3994 7030 -3960
rect 6833 -4011 7030 -3994
rect -1110 -4028 7030 -4011
rect -1110 -4030 -1070 -4028
rect -1104 -4062 -1070 -4030
rect -1036 -4030 -428 -4028
rect -1036 -4062 -1003 -4030
rect -1104 -4262 -1003 -4062
rect -1104 -4296 -1070 -4262
rect -1036 -4296 -1003 -4262
rect -1104 -4330 -1003 -4296
rect -1104 -4364 -1070 -4330
rect -1036 -4364 -1003 -4330
rect -1104 -4398 -1003 -4364
rect -941 -4045 -869 -4030
rect -941 -4079 -917 -4045
rect -883 -4079 -869 -4045
rect -941 -4245 -869 -4079
rect -595 -4045 -523 -4030
rect -595 -4079 -581 -4045
rect -547 -4079 -523 -4045
rect -811 -4097 -653 -4083
rect -811 -4131 -797 -4097
rect -763 -4111 -701 -4097
rect -667 -4131 -653 -4097
rect -811 -4193 -783 -4131
rect -681 -4193 -653 -4131
rect -811 -4227 -797 -4193
rect -763 -4227 -701 -4213
rect -667 -4227 -653 -4193
rect -811 -4241 -653 -4227
rect -941 -4279 -917 -4245
rect -883 -4279 -869 -4245
rect -941 -4299 -869 -4279
rect -595 -4245 -523 -4079
rect -595 -4279 -581 -4245
rect -547 -4279 -523 -4245
rect -595 -4299 -523 -4279
rect -941 -4313 -523 -4299
rect -941 -4347 -917 -4313
rect -883 -4347 -849 -4313
rect -815 -4347 -649 -4313
rect -615 -4347 -581 -4313
rect -547 -4347 -523 -4313
rect -941 -4371 -523 -4347
rect -461 -4062 -428 -4030
rect -394 -4030 -250 -4028
rect -394 -4062 -360 -4030
rect -461 -4262 -360 -4062
rect -461 -4296 -428 -4262
rect -394 -4296 -360 -4262
rect -461 -4330 -360 -4296
rect -461 -4364 -428 -4330
rect -394 -4364 -360 -4330
rect -1104 -4432 -1070 -4398
rect -1036 -4432 -1003 -4398
rect -1104 -4433 -1003 -4432
rect -461 -4398 -360 -4364
rect -461 -4432 -428 -4398
rect -394 -4432 -360 -4398
rect -461 -4433 -360 -4432
rect -1104 -4466 -360 -4433
rect -1104 -4500 -1070 -4466
rect -1036 -4500 -1002 -4466
rect -968 -4500 -934 -4466
rect -900 -4500 -866 -4466
rect -832 -4500 -632 -4466
rect -598 -4500 -564 -4466
rect -530 -4500 -496 -4466
rect -462 -4500 -428 -4466
rect -394 -4500 -360 -4466
rect -1104 -4534 -360 -4500
rect -284 -4062 -250 -4030
rect -216 -4030 392 -4028
rect -216 -4062 -183 -4030
rect -284 -4262 -183 -4062
rect -284 -4296 -250 -4262
rect -216 -4296 -183 -4262
rect -284 -4330 -183 -4296
rect -284 -4364 -250 -4330
rect -216 -4364 -183 -4330
rect -284 -4398 -183 -4364
rect -121 -4045 -49 -4030
rect -121 -4079 -97 -4045
rect -63 -4079 -49 -4045
rect -121 -4245 -49 -4079
rect 225 -4045 297 -4030
rect 225 -4079 239 -4045
rect 273 -4079 297 -4045
rect 9 -4097 167 -4083
rect 9 -4131 23 -4097
rect 57 -4111 119 -4097
rect 153 -4131 167 -4097
rect 9 -4193 37 -4131
rect 139 -4193 167 -4131
rect 9 -4227 23 -4193
rect 57 -4227 119 -4213
rect 153 -4227 167 -4193
rect 9 -4241 167 -4227
rect -121 -4279 -97 -4245
rect -63 -4279 -49 -4245
rect -121 -4299 -49 -4279
rect 225 -4245 297 -4079
rect 225 -4279 239 -4245
rect 273 -4279 297 -4245
rect 225 -4299 297 -4279
rect -121 -4313 297 -4299
rect -121 -4347 -97 -4313
rect -63 -4347 -29 -4313
rect 5 -4347 171 -4313
rect 205 -4347 239 -4313
rect 273 -4347 297 -4313
rect -121 -4371 297 -4347
rect 359 -4062 392 -4030
rect 426 -4030 570 -4028
rect 426 -4062 460 -4030
rect 359 -4262 460 -4062
rect 359 -4296 392 -4262
rect 426 -4296 460 -4262
rect 359 -4330 460 -4296
rect 359 -4364 392 -4330
rect 426 -4364 460 -4330
rect -284 -4432 -250 -4398
rect -216 -4432 -183 -4398
rect -284 -4433 -183 -4432
rect 359 -4398 460 -4364
rect 359 -4432 392 -4398
rect 426 -4432 460 -4398
rect 359 -4433 460 -4432
rect -284 -4466 460 -4433
rect -284 -4500 -250 -4466
rect -216 -4500 -182 -4466
rect -148 -4500 -114 -4466
rect -80 -4500 -46 -4466
rect -12 -4500 188 -4466
rect 222 -4500 256 -4466
rect 290 -4500 324 -4466
rect 358 -4500 392 -4466
rect 426 -4500 460 -4466
rect -284 -4534 460 -4500
rect 536 -4062 570 -4030
rect 604 -4030 1212 -4028
rect 604 -4062 637 -4030
rect 536 -4262 637 -4062
rect 536 -4296 570 -4262
rect 604 -4296 637 -4262
rect 536 -4330 637 -4296
rect 536 -4364 570 -4330
rect 604 -4364 637 -4330
rect 536 -4398 637 -4364
rect 699 -4045 771 -4030
rect 699 -4079 723 -4045
rect 757 -4079 771 -4045
rect 699 -4245 771 -4079
rect 1045 -4045 1117 -4030
rect 1045 -4079 1059 -4045
rect 1093 -4079 1117 -4045
rect 829 -4097 987 -4083
rect 829 -4131 843 -4097
rect 877 -4111 939 -4097
rect 973 -4131 987 -4097
rect 829 -4193 857 -4131
rect 959 -4193 987 -4131
rect 829 -4227 843 -4193
rect 877 -4227 939 -4213
rect 973 -4227 987 -4193
rect 829 -4241 987 -4227
rect 699 -4279 723 -4245
rect 757 -4279 771 -4245
rect 699 -4299 771 -4279
rect 1045 -4245 1117 -4079
rect 1045 -4279 1059 -4245
rect 1093 -4279 1117 -4245
rect 1045 -4299 1117 -4279
rect 699 -4313 1117 -4299
rect 699 -4347 723 -4313
rect 757 -4347 791 -4313
rect 825 -4347 991 -4313
rect 1025 -4347 1059 -4313
rect 1093 -4347 1117 -4313
rect 699 -4371 1117 -4347
rect 1179 -4062 1212 -4030
rect 1246 -4030 1390 -4028
rect 1246 -4062 1280 -4030
rect 1179 -4262 1280 -4062
rect 1179 -4296 1212 -4262
rect 1246 -4296 1280 -4262
rect 1179 -4330 1280 -4296
rect 1179 -4364 1212 -4330
rect 1246 -4364 1280 -4330
rect 536 -4432 570 -4398
rect 604 -4432 637 -4398
rect 536 -4433 637 -4432
rect 1179 -4398 1280 -4364
rect 1179 -4432 1212 -4398
rect 1246 -4432 1280 -4398
rect 1179 -4433 1280 -4432
rect 536 -4466 1280 -4433
rect 536 -4500 570 -4466
rect 604 -4500 638 -4466
rect 672 -4500 706 -4466
rect 740 -4500 774 -4466
rect 808 -4500 1008 -4466
rect 1042 -4500 1076 -4466
rect 1110 -4500 1144 -4466
rect 1178 -4500 1212 -4466
rect 1246 -4500 1280 -4466
rect 536 -4534 1280 -4500
rect 1356 -4062 1390 -4030
rect 1424 -4030 2032 -4028
rect 1424 -4062 1457 -4030
rect 1356 -4262 1457 -4062
rect 1356 -4296 1390 -4262
rect 1424 -4296 1457 -4262
rect 1356 -4330 1457 -4296
rect 1356 -4364 1390 -4330
rect 1424 -4364 1457 -4330
rect 1356 -4398 1457 -4364
rect 1519 -4045 1591 -4030
rect 1519 -4079 1543 -4045
rect 1577 -4079 1591 -4045
rect 1519 -4245 1591 -4079
rect 1865 -4045 1937 -4030
rect 1865 -4079 1879 -4045
rect 1913 -4079 1937 -4045
rect 1649 -4097 1807 -4083
rect 1649 -4131 1663 -4097
rect 1697 -4111 1759 -4097
rect 1793 -4131 1807 -4097
rect 1649 -4193 1677 -4131
rect 1779 -4193 1807 -4131
rect 1649 -4227 1663 -4193
rect 1697 -4227 1759 -4213
rect 1793 -4227 1807 -4193
rect 1649 -4241 1807 -4227
rect 1519 -4279 1543 -4245
rect 1577 -4279 1591 -4245
rect 1519 -4299 1591 -4279
rect 1865 -4245 1937 -4079
rect 1865 -4279 1879 -4245
rect 1913 -4279 1937 -4245
rect 1865 -4299 1937 -4279
rect 1519 -4313 1937 -4299
rect 1519 -4347 1543 -4313
rect 1577 -4347 1611 -4313
rect 1645 -4347 1811 -4313
rect 1845 -4347 1879 -4313
rect 1913 -4347 1937 -4313
rect 1519 -4371 1937 -4347
rect 1999 -4062 2032 -4030
rect 2066 -4030 2210 -4028
rect 2066 -4062 2100 -4030
rect 1999 -4262 2100 -4062
rect 1999 -4296 2032 -4262
rect 2066 -4296 2100 -4262
rect 1999 -4330 2100 -4296
rect 1999 -4364 2032 -4330
rect 2066 -4364 2100 -4330
rect 1356 -4432 1390 -4398
rect 1424 -4432 1457 -4398
rect 1356 -4433 1457 -4432
rect 1999 -4398 2100 -4364
rect 1999 -4432 2032 -4398
rect 2066 -4432 2100 -4398
rect 1999 -4433 2100 -4432
rect 1356 -4466 2100 -4433
rect 1356 -4500 1390 -4466
rect 1424 -4500 1458 -4466
rect 1492 -4500 1526 -4466
rect 1560 -4500 1594 -4466
rect 1628 -4500 1828 -4466
rect 1862 -4500 1896 -4466
rect 1930 -4500 1964 -4466
rect 1998 -4500 2032 -4466
rect 2066 -4500 2100 -4466
rect 1356 -4534 2100 -4500
rect 2176 -4062 2210 -4030
rect 2244 -4030 2852 -4028
rect 2244 -4062 2277 -4030
rect 2176 -4262 2277 -4062
rect 2176 -4296 2210 -4262
rect 2244 -4296 2277 -4262
rect 2176 -4330 2277 -4296
rect 2176 -4364 2210 -4330
rect 2244 -4364 2277 -4330
rect 2176 -4398 2277 -4364
rect 2339 -4045 2411 -4030
rect 2339 -4079 2363 -4045
rect 2397 -4079 2411 -4045
rect 2339 -4245 2411 -4079
rect 2685 -4045 2757 -4030
rect 2685 -4079 2699 -4045
rect 2733 -4079 2757 -4045
rect 2469 -4097 2627 -4083
rect 2469 -4131 2483 -4097
rect 2517 -4111 2579 -4097
rect 2613 -4131 2627 -4097
rect 2469 -4193 2497 -4131
rect 2599 -4193 2627 -4131
rect 2469 -4227 2483 -4193
rect 2517 -4227 2579 -4213
rect 2613 -4227 2627 -4193
rect 2469 -4241 2627 -4227
rect 2339 -4279 2363 -4245
rect 2397 -4279 2411 -4245
rect 2339 -4299 2411 -4279
rect 2685 -4245 2757 -4079
rect 2685 -4279 2699 -4245
rect 2733 -4279 2757 -4245
rect 2685 -4299 2757 -4279
rect 2339 -4313 2757 -4299
rect 2339 -4347 2363 -4313
rect 2397 -4347 2431 -4313
rect 2465 -4347 2631 -4313
rect 2665 -4347 2699 -4313
rect 2733 -4347 2757 -4313
rect 2339 -4371 2757 -4347
rect 2819 -4062 2852 -4030
rect 2886 -4030 3030 -4028
rect 2886 -4062 2920 -4030
rect 2819 -4262 2920 -4062
rect 2819 -4296 2852 -4262
rect 2886 -4296 2920 -4262
rect 2819 -4330 2920 -4296
rect 2819 -4364 2852 -4330
rect 2886 -4364 2920 -4330
rect 2176 -4432 2210 -4398
rect 2244 -4432 2277 -4398
rect 2176 -4433 2277 -4432
rect 2819 -4398 2920 -4364
rect 2819 -4432 2852 -4398
rect 2886 -4432 2920 -4398
rect 2819 -4433 2920 -4432
rect 2176 -4466 2920 -4433
rect 2176 -4500 2210 -4466
rect 2244 -4500 2278 -4466
rect 2312 -4500 2346 -4466
rect 2380 -4500 2414 -4466
rect 2448 -4500 2648 -4466
rect 2682 -4500 2716 -4466
rect 2750 -4500 2784 -4466
rect 2818 -4500 2852 -4466
rect 2886 -4500 2920 -4466
rect 2176 -4534 2920 -4500
rect 2996 -4062 3030 -4030
rect 3064 -4030 3672 -4028
rect 3064 -4062 3097 -4030
rect 2996 -4262 3097 -4062
rect 2996 -4296 3030 -4262
rect 3064 -4296 3097 -4262
rect 2996 -4330 3097 -4296
rect 2996 -4364 3030 -4330
rect 3064 -4364 3097 -4330
rect 2996 -4398 3097 -4364
rect 3159 -4045 3231 -4030
rect 3159 -4079 3183 -4045
rect 3217 -4079 3231 -4045
rect 3159 -4245 3231 -4079
rect 3505 -4045 3577 -4030
rect 3505 -4079 3519 -4045
rect 3553 -4079 3577 -4045
rect 3289 -4097 3447 -4083
rect 3289 -4131 3303 -4097
rect 3337 -4111 3399 -4097
rect 3433 -4131 3447 -4097
rect 3289 -4193 3317 -4131
rect 3419 -4193 3447 -4131
rect 3289 -4227 3303 -4193
rect 3337 -4227 3399 -4213
rect 3433 -4227 3447 -4193
rect 3289 -4241 3447 -4227
rect 3159 -4279 3183 -4245
rect 3217 -4279 3231 -4245
rect 3159 -4299 3231 -4279
rect 3505 -4245 3577 -4079
rect 3505 -4279 3519 -4245
rect 3553 -4279 3577 -4245
rect 3505 -4299 3577 -4279
rect 3159 -4313 3577 -4299
rect 3159 -4347 3183 -4313
rect 3217 -4347 3251 -4313
rect 3285 -4347 3451 -4313
rect 3485 -4347 3519 -4313
rect 3553 -4347 3577 -4313
rect 3159 -4371 3577 -4347
rect 3639 -4062 3672 -4030
rect 3706 -4030 3850 -4028
rect 3706 -4062 3740 -4030
rect 3639 -4262 3740 -4062
rect 3639 -4296 3672 -4262
rect 3706 -4296 3740 -4262
rect 3639 -4330 3740 -4296
rect 3639 -4364 3672 -4330
rect 3706 -4364 3740 -4330
rect 2996 -4432 3030 -4398
rect 3064 -4432 3097 -4398
rect 2996 -4433 3097 -4432
rect 3639 -4398 3740 -4364
rect 3639 -4432 3672 -4398
rect 3706 -4432 3740 -4398
rect 3639 -4433 3740 -4432
rect 2996 -4466 3740 -4433
rect 2996 -4500 3030 -4466
rect 3064 -4500 3098 -4466
rect 3132 -4500 3166 -4466
rect 3200 -4500 3234 -4466
rect 3268 -4500 3468 -4466
rect 3502 -4500 3536 -4466
rect 3570 -4500 3604 -4466
rect 3638 -4500 3672 -4466
rect 3706 -4500 3740 -4466
rect 2996 -4534 3740 -4500
rect 3816 -4062 3850 -4030
rect 3884 -4030 4492 -4028
rect 3884 -4062 3917 -4030
rect 3816 -4262 3917 -4062
rect 3816 -4296 3850 -4262
rect 3884 -4296 3917 -4262
rect 3816 -4330 3917 -4296
rect 3816 -4364 3850 -4330
rect 3884 -4364 3917 -4330
rect 3816 -4398 3917 -4364
rect 3979 -4045 4051 -4030
rect 3979 -4079 4003 -4045
rect 4037 -4079 4051 -4045
rect 3979 -4245 4051 -4079
rect 4325 -4045 4397 -4030
rect 4325 -4079 4339 -4045
rect 4373 -4079 4397 -4045
rect 4109 -4097 4267 -4083
rect 4109 -4131 4123 -4097
rect 4157 -4111 4219 -4097
rect 4253 -4131 4267 -4097
rect 4109 -4193 4137 -4131
rect 4239 -4193 4267 -4131
rect 4109 -4227 4123 -4193
rect 4157 -4227 4219 -4213
rect 4253 -4227 4267 -4193
rect 4109 -4241 4267 -4227
rect 3979 -4279 4003 -4245
rect 4037 -4279 4051 -4245
rect 3979 -4299 4051 -4279
rect 4325 -4245 4397 -4079
rect 4325 -4279 4339 -4245
rect 4373 -4279 4397 -4245
rect 4325 -4299 4397 -4279
rect 3979 -4313 4397 -4299
rect 3979 -4347 4003 -4313
rect 4037 -4347 4071 -4313
rect 4105 -4347 4271 -4313
rect 4305 -4347 4339 -4313
rect 4373 -4347 4397 -4313
rect 3979 -4371 4397 -4347
rect 4459 -4062 4492 -4030
rect 4526 -4030 4670 -4028
rect 4526 -4062 4560 -4030
rect 4459 -4262 4560 -4062
rect 4459 -4296 4492 -4262
rect 4526 -4296 4560 -4262
rect 4459 -4330 4560 -4296
rect 4459 -4364 4492 -4330
rect 4526 -4364 4560 -4330
rect 3816 -4432 3850 -4398
rect 3884 -4432 3917 -4398
rect 3816 -4433 3917 -4432
rect 4459 -4398 4560 -4364
rect 4459 -4432 4492 -4398
rect 4526 -4432 4560 -4398
rect 4459 -4433 4560 -4432
rect 3816 -4466 4560 -4433
rect 3816 -4500 3850 -4466
rect 3884 -4500 3918 -4466
rect 3952 -4500 3986 -4466
rect 4020 -4500 4054 -4466
rect 4088 -4500 4288 -4466
rect 4322 -4500 4356 -4466
rect 4390 -4500 4424 -4466
rect 4458 -4500 4492 -4466
rect 4526 -4500 4560 -4466
rect 3816 -4534 4560 -4500
rect 4636 -4062 4670 -4030
rect 4704 -4030 5312 -4028
rect 4704 -4062 4737 -4030
rect 4636 -4262 4737 -4062
rect 4636 -4296 4670 -4262
rect 4704 -4296 4737 -4262
rect 4636 -4330 4737 -4296
rect 4636 -4364 4670 -4330
rect 4704 -4364 4737 -4330
rect 4636 -4398 4737 -4364
rect 4799 -4045 4871 -4030
rect 4799 -4079 4823 -4045
rect 4857 -4079 4871 -4045
rect 4799 -4245 4871 -4079
rect 5145 -4045 5217 -4030
rect 5145 -4079 5159 -4045
rect 5193 -4079 5217 -4045
rect 4929 -4097 5087 -4083
rect 4929 -4131 4943 -4097
rect 4977 -4111 5039 -4097
rect 5073 -4131 5087 -4097
rect 4929 -4193 4957 -4131
rect 5059 -4193 5087 -4131
rect 4929 -4227 4943 -4193
rect 4977 -4227 5039 -4213
rect 5073 -4227 5087 -4193
rect 4929 -4241 5087 -4227
rect 4799 -4279 4823 -4245
rect 4857 -4279 4871 -4245
rect 4799 -4299 4871 -4279
rect 5145 -4245 5217 -4079
rect 5145 -4279 5159 -4245
rect 5193 -4279 5217 -4245
rect 5145 -4299 5217 -4279
rect 4799 -4313 5217 -4299
rect 4799 -4347 4823 -4313
rect 4857 -4347 4891 -4313
rect 4925 -4347 5091 -4313
rect 5125 -4347 5159 -4313
rect 5193 -4347 5217 -4313
rect 4799 -4371 5217 -4347
rect 5279 -4062 5312 -4030
rect 5346 -4030 5490 -4028
rect 5346 -4062 5380 -4030
rect 5279 -4262 5380 -4062
rect 5279 -4296 5312 -4262
rect 5346 -4296 5380 -4262
rect 5279 -4330 5380 -4296
rect 5279 -4364 5312 -4330
rect 5346 -4364 5380 -4330
rect 4636 -4432 4670 -4398
rect 4704 -4432 4737 -4398
rect 4636 -4433 4737 -4432
rect 5279 -4398 5380 -4364
rect 5279 -4432 5312 -4398
rect 5346 -4432 5380 -4398
rect 5279 -4433 5380 -4432
rect 4636 -4466 5380 -4433
rect 4636 -4500 4670 -4466
rect 4704 -4500 4738 -4466
rect 4772 -4500 4806 -4466
rect 4840 -4500 4874 -4466
rect 4908 -4500 5108 -4466
rect 5142 -4500 5176 -4466
rect 5210 -4500 5244 -4466
rect 5278 -4500 5312 -4466
rect 5346 -4500 5380 -4466
rect 4636 -4534 5380 -4500
rect 5456 -4062 5490 -4030
rect 5524 -4030 6132 -4028
rect 5524 -4062 5557 -4030
rect 5456 -4262 5557 -4062
rect 5456 -4296 5490 -4262
rect 5524 -4296 5557 -4262
rect 5456 -4330 5557 -4296
rect 5456 -4364 5490 -4330
rect 5524 -4364 5557 -4330
rect 5456 -4398 5557 -4364
rect 5619 -4045 5691 -4030
rect 5619 -4079 5643 -4045
rect 5677 -4079 5691 -4045
rect 5619 -4245 5691 -4079
rect 5965 -4045 6037 -4030
rect 5965 -4079 5979 -4045
rect 6013 -4079 6037 -4045
rect 5749 -4097 5907 -4083
rect 5749 -4131 5763 -4097
rect 5797 -4111 5859 -4097
rect 5893 -4131 5907 -4097
rect 5749 -4193 5777 -4131
rect 5879 -4193 5907 -4131
rect 5749 -4227 5763 -4193
rect 5797 -4227 5859 -4213
rect 5893 -4227 5907 -4193
rect 5749 -4241 5907 -4227
rect 5619 -4279 5643 -4245
rect 5677 -4279 5691 -4245
rect 5619 -4299 5691 -4279
rect 5965 -4245 6037 -4079
rect 5965 -4279 5979 -4245
rect 6013 -4279 6037 -4245
rect 5965 -4299 6037 -4279
rect 5619 -4313 6037 -4299
rect 5619 -4347 5643 -4313
rect 5677 -4347 5711 -4313
rect 5745 -4347 5911 -4313
rect 5945 -4347 5979 -4313
rect 6013 -4347 6037 -4313
rect 5619 -4371 6037 -4347
rect 6099 -4062 6132 -4030
rect 6166 -4030 6310 -4028
rect 6166 -4062 6200 -4030
rect 6099 -4262 6200 -4062
rect 6099 -4296 6132 -4262
rect 6166 -4296 6200 -4262
rect 6099 -4330 6200 -4296
rect 6099 -4364 6132 -4330
rect 6166 -4364 6200 -4330
rect 5456 -4432 5490 -4398
rect 5524 -4432 5557 -4398
rect 5456 -4433 5557 -4432
rect 6099 -4398 6200 -4364
rect 6099 -4432 6132 -4398
rect 6166 -4432 6200 -4398
rect 6099 -4433 6200 -4432
rect 5456 -4466 6200 -4433
rect 5456 -4500 5490 -4466
rect 5524 -4500 5558 -4466
rect 5592 -4500 5626 -4466
rect 5660 -4500 5694 -4466
rect 5728 -4500 5928 -4466
rect 5962 -4500 5996 -4466
rect 6030 -4500 6064 -4466
rect 6098 -4500 6132 -4466
rect 6166 -4500 6200 -4466
rect 5456 -4534 6200 -4500
rect 6276 -4062 6310 -4030
rect 6344 -4030 6952 -4028
rect 6344 -4062 6377 -4030
rect 6276 -4262 6377 -4062
rect 6276 -4296 6310 -4262
rect 6344 -4296 6377 -4262
rect 6276 -4330 6377 -4296
rect 6276 -4364 6310 -4330
rect 6344 -4364 6377 -4330
rect 6276 -4398 6377 -4364
rect 6439 -4045 6511 -4030
rect 6439 -4079 6463 -4045
rect 6497 -4079 6511 -4045
rect 6439 -4245 6511 -4079
rect 6785 -4045 6857 -4030
rect 6785 -4079 6799 -4045
rect 6833 -4079 6857 -4045
rect 6569 -4097 6727 -4083
rect 6569 -4131 6583 -4097
rect 6617 -4111 6679 -4097
rect 6713 -4131 6727 -4097
rect 6569 -4193 6597 -4131
rect 6699 -4193 6727 -4131
rect 6569 -4227 6583 -4193
rect 6617 -4227 6679 -4213
rect 6713 -4227 6727 -4193
rect 6569 -4241 6727 -4227
rect 6439 -4279 6463 -4245
rect 6497 -4279 6511 -4245
rect 6439 -4299 6511 -4279
rect 6785 -4245 6857 -4079
rect 6785 -4279 6799 -4245
rect 6833 -4279 6857 -4245
rect 6785 -4299 6857 -4279
rect 6439 -4313 6857 -4299
rect 6439 -4347 6463 -4313
rect 6497 -4347 6531 -4313
rect 6565 -4347 6731 -4313
rect 6765 -4347 6799 -4313
rect 6833 -4347 6857 -4313
rect 6439 -4371 6857 -4347
rect 6919 -4062 6952 -4030
rect 6986 -4030 7030 -4028
rect 6986 -4062 7020 -4030
rect 6919 -4262 7020 -4062
rect 6919 -4296 6952 -4262
rect 6986 -4296 7020 -4262
rect 6919 -4330 7020 -4296
rect 6919 -4364 6952 -4330
rect 6986 -4364 7020 -4330
rect 6276 -4432 6310 -4398
rect 6344 -4432 6377 -4398
rect 6276 -4433 6377 -4432
rect 6919 -4398 7020 -4364
rect 6919 -4432 6952 -4398
rect 6986 -4432 7020 -4398
rect 6919 -4433 7020 -4432
rect 6276 -4466 7020 -4433
rect 6276 -4500 6310 -4466
rect 6344 -4500 6378 -4466
rect 6412 -4500 6446 -4466
rect 6480 -4500 6514 -4466
rect 6548 -4500 6748 -4466
rect 6782 -4500 6816 -4466
rect 6850 -4500 6884 -4466
rect 6918 -4500 6952 -4466
rect 6986 -4500 7020 -4466
rect 6276 -4534 7020 -4500
rect 15760 -4810 15840 -3320
<< viali >>
rect 6720 4360 6760 4400
rect 7560 4300 7600 6240
rect 7660 4300 7700 6240
rect 7760 4300 7800 6240
rect 8070 4650 8110 4690
rect 7500 4150 7540 4190
rect 7820 4150 7860 4190
rect 7260 3920 7300 3960
rect 7560 2090 7600 4030
rect 7660 2090 7700 4030
rect 7760 2090 7800 4030
rect 8650 2830 8730 2910
rect 12110 2830 12490 2910
rect 15740 2830 16120 2910
rect 17030 2830 17410 2910
rect 15880 1220 15920 1260
rect 15850 780 15920 930
rect 7260 570 7300 610
rect 7670 570 7710 610
rect 6650 40 6730 420
rect 7850 40 7930 420
rect -797 -831 -763 -817
rect -701 -831 -667 -817
rect -797 -851 -783 -831
rect -783 -851 -763 -831
rect -701 -851 -681 -831
rect -681 -851 -667 -831
rect -797 -933 -783 -913
rect -783 -933 -763 -913
rect -701 -933 -681 -913
rect -681 -933 -667 -913
rect -797 -947 -763 -933
rect -701 -947 -667 -933
rect 23 -831 57 -817
rect 119 -831 153 -817
rect 23 -851 37 -831
rect 37 -851 57 -831
rect 119 -851 139 -831
rect 139 -851 153 -831
rect 23 -933 37 -913
rect 37 -933 57 -913
rect 119 -933 139 -913
rect 139 -933 153 -913
rect 23 -947 57 -933
rect 119 -947 153 -933
rect 843 -831 877 -817
rect 939 -831 973 -817
rect 843 -851 857 -831
rect 857 -851 877 -831
rect 939 -851 959 -831
rect 959 -851 973 -831
rect 843 -933 857 -913
rect 857 -933 877 -913
rect 939 -933 959 -913
rect 959 -933 973 -913
rect 843 -947 877 -933
rect 939 -947 973 -933
rect 1663 -831 1697 -817
rect 1759 -831 1793 -817
rect 1663 -851 1677 -831
rect 1677 -851 1697 -831
rect 1759 -851 1779 -831
rect 1779 -851 1793 -831
rect 1663 -933 1677 -913
rect 1677 -933 1697 -913
rect 1759 -933 1779 -913
rect 1779 -933 1793 -913
rect 1663 -947 1697 -933
rect 1759 -947 1793 -933
rect 2483 -831 2517 -817
rect 2579 -831 2613 -817
rect 2483 -851 2497 -831
rect 2497 -851 2517 -831
rect 2579 -851 2599 -831
rect 2599 -851 2613 -831
rect 2483 -933 2497 -913
rect 2497 -933 2517 -913
rect 2579 -933 2599 -913
rect 2599 -933 2613 -913
rect 2483 -947 2517 -933
rect 2579 -947 2613 -933
rect 3303 -831 3337 -817
rect 3399 -831 3433 -817
rect 3303 -851 3317 -831
rect 3317 -851 3337 -831
rect 3399 -851 3419 -831
rect 3419 -851 3433 -831
rect 3303 -933 3317 -913
rect 3317 -933 3337 -913
rect 3399 -933 3419 -913
rect 3419 -933 3433 -913
rect 3303 -947 3337 -933
rect 3399 -947 3433 -933
rect 4123 -831 4157 -817
rect 4219 -831 4253 -817
rect 4123 -851 4137 -831
rect 4137 -851 4157 -831
rect 4219 -851 4239 -831
rect 4239 -851 4253 -831
rect 4123 -933 4137 -913
rect 4137 -933 4157 -913
rect 4219 -933 4239 -913
rect 4239 -933 4253 -913
rect 4123 -947 4157 -933
rect 4219 -947 4253 -933
rect 4943 -831 4977 -817
rect 5039 -831 5073 -817
rect 4943 -851 4957 -831
rect 4957 -851 4977 -831
rect 5039 -851 5059 -831
rect 5059 -851 5073 -831
rect 4943 -933 4957 -913
rect 4957 -933 4977 -913
rect 5039 -933 5059 -913
rect 5059 -933 5073 -913
rect 4943 -947 4977 -933
rect 5039 -947 5073 -933
rect 5763 -831 5797 -817
rect 5859 -831 5893 -817
rect 5763 -851 5777 -831
rect 5777 -851 5797 -831
rect 5859 -851 5879 -831
rect 5879 -851 5893 -831
rect 5763 -933 5777 -913
rect 5777 -933 5797 -913
rect 5859 -933 5879 -913
rect 5879 -933 5893 -913
rect 5763 -947 5797 -933
rect 5859 -947 5893 -933
rect 6583 -831 6617 -817
rect 6679 -831 6713 -817
rect 6583 -851 6597 -831
rect 6597 -851 6617 -831
rect 6679 -851 6699 -831
rect 6699 -851 6713 -831
rect 6583 -933 6597 -913
rect 6597 -933 6617 -913
rect 6679 -933 6699 -913
rect 6699 -933 6713 -913
rect 6583 -947 6617 -933
rect 6679 -947 6713 -933
rect 7433 -831 7467 -817
rect 7529 -831 7563 -817
rect 7433 -851 7447 -831
rect 7447 -851 7467 -831
rect 7529 -851 7549 -831
rect 7549 -851 7563 -831
rect 7433 -933 7447 -913
rect 7447 -933 7467 -913
rect 7529 -933 7549 -913
rect 7549 -933 7563 -913
rect 7433 -947 7467 -933
rect 7529 -947 7563 -933
rect -797 -1651 -763 -1637
rect -701 -1651 -667 -1637
rect -797 -1671 -783 -1651
rect -783 -1671 -763 -1651
rect -701 -1671 -681 -1651
rect -681 -1671 -667 -1651
rect -797 -1753 -783 -1733
rect -783 -1753 -763 -1733
rect -701 -1753 -681 -1733
rect -681 -1753 -667 -1733
rect -797 -1767 -763 -1753
rect -701 -1767 -667 -1753
rect 23 -1651 57 -1637
rect 119 -1651 153 -1637
rect 23 -1671 37 -1651
rect 37 -1671 57 -1651
rect 119 -1671 139 -1651
rect 139 -1671 153 -1651
rect 23 -1753 37 -1733
rect 37 -1753 57 -1733
rect 119 -1753 139 -1733
rect 139 -1753 153 -1733
rect 23 -1767 57 -1753
rect 119 -1767 153 -1753
rect 843 -1651 877 -1637
rect 939 -1651 973 -1637
rect 843 -1671 857 -1651
rect 857 -1671 877 -1651
rect 939 -1671 959 -1651
rect 959 -1671 973 -1651
rect 843 -1753 857 -1733
rect 857 -1753 877 -1733
rect 939 -1753 959 -1733
rect 959 -1753 973 -1733
rect 843 -1767 877 -1753
rect 939 -1767 973 -1753
rect 1663 -1651 1697 -1637
rect 1759 -1651 1793 -1637
rect 1663 -1671 1677 -1651
rect 1677 -1671 1697 -1651
rect 1759 -1671 1779 -1651
rect 1779 -1671 1793 -1651
rect 1663 -1753 1677 -1733
rect 1677 -1753 1697 -1733
rect 1759 -1753 1779 -1733
rect 1779 -1753 1793 -1733
rect 1663 -1767 1697 -1753
rect 1759 -1767 1793 -1753
rect 2483 -1651 2517 -1637
rect 2579 -1651 2613 -1637
rect 2483 -1671 2497 -1651
rect 2497 -1671 2517 -1651
rect 2579 -1671 2599 -1651
rect 2599 -1671 2613 -1651
rect 2483 -1753 2497 -1733
rect 2497 -1753 2517 -1733
rect 2579 -1753 2599 -1733
rect 2599 -1753 2613 -1733
rect 2483 -1767 2517 -1753
rect 2579 -1767 2613 -1753
rect 3303 -1651 3337 -1637
rect 3399 -1651 3433 -1637
rect 3303 -1671 3317 -1651
rect 3317 -1671 3337 -1651
rect 3399 -1671 3419 -1651
rect 3419 -1671 3433 -1651
rect 3303 -1753 3317 -1733
rect 3317 -1753 3337 -1733
rect 3399 -1753 3419 -1733
rect 3419 -1753 3433 -1733
rect 3303 -1767 3337 -1753
rect 3399 -1767 3433 -1753
rect 4123 -1651 4157 -1637
rect 4219 -1651 4253 -1637
rect 4123 -1671 4137 -1651
rect 4137 -1671 4157 -1651
rect 4219 -1671 4239 -1651
rect 4239 -1671 4253 -1651
rect 4123 -1753 4137 -1733
rect 4137 -1753 4157 -1733
rect 4219 -1753 4239 -1733
rect 4239 -1753 4253 -1733
rect 4123 -1767 4157 -1753
rect 4219 -1767 4253 -1753
rect 4943 -1651 4977 -1637
rect 5039 -1651 5073 -1637
rect 4943 -1671 4957 -1651
rect 4957 -1671 4977 -1651
rect 5039 -1671 5059 -1651
rect 5059 -1671 5073 -1651
rect 4943 -1753 4957 -1733
rect 4957 -1753 4977 -1733
rect 5039 -1753 5059 -1733
rect 5059 -1753 5073 -1733
rect 4943 -1767 4977 -1753
rect 5039 -1767 5073 -1753
rect 5763 -1651 5797 -1637
rect 5859 -1651 5893 -1637
rect 5763 -1671 5777 -1651
rect 5777 -1671 5797 -1651
rect 5859 -1671 5879 -1651
rect 5879 -1671 5893 -1651
rect 5763 -1753 5777 -1733
rect 5777 -1753 5797 -1733
rect 5859 -1753 5879 -1733
rect 5879 -1753 5893 -1733
rect 5763 -1767 5797 -1753
rect 5859 -1767 5893 -1753
rect 6583 -1651 6617 -1637
rect 6679 -1651 6713 -1637
rect 6583 -1671 6597 -1651
rect 6597 -1671 6617 -1651
rect 6679 -1671 6699 -1651
rect 6699 -1671 6713 -1651
rect 6583 -1753 6597 -1733
rect 6597 -1753 6617 -1733
rect 6679 -1753 6699 -1733
rect 6699 -1753 6713 -1733
rect 6583 -1767 6617 -1753
rect 6679 -1767 6713 -1753
rect 8620 -1630 8760 -1170
rect 17000 -1310 17080 -930
rect -797 -2471 -763 -2457
rect -701 -2471 -667 -2457
rect -797 -2491 -783 -2471
rect -783 -2491 -763 -2471
rect -701 -2491 -681 -2471
rect -681 -2491 -667 -2471
rect -797 -2573 -783 -2553
rect -783 -2573 -763 -2553
rect -701 -2573 -681 -2553
rect -681 -2573 -667 -2553
rect -797 -2587 -763 -2573
rect -701 -2587 -667 -2573
rect 23 -2471 57 -2457
rect 119 -2471 153 -2457
rect 23 -2491 37 -2471
rect 37 -2491 57 -2471
rect 119 -2491 139 -2471
rect 139 -2491 153 -2471
rect 23 -2573 37 -2553
rect 37 -2573 57 -2553
rect 119 -2573 139 -2553
rect 139 -2573 153 -2553
rect 23 -2587 57 -2573
rect 119 -2587 153 -2573
rect 843 -2471 877 -2457
rect 939 -2471 973 -2457
rect 843 -2491 857 -2471
rect 857 -2491 877 -2471
rect 939 -2491 959 -2471
rect 959 -2491 973 -2471
rect 843 -2573 857 -2553
rect 857 -2573 877 -2553
rect 939 -2573 959 -2553
rect 959 -2573 973 -2553
rect 843 -2587 877 -2573
rect 939 -2587 973 -2573
rect 1663 -2471 1697 -2457
rect 1759 -2471 1793 -2457
rect 1663 -2491 1677 -2471
rect 1677 -2491 1697 -2471
rect 1759 -2491 1779 -2471
rect 1779 -2491 1793 -2471
rect 1663 -2573 1677 -2553
rect 1677 -2573 1697 -2553
rect 1759 -2573 1779 -2553
rect 1779 -2573 1793 -2553
rect 1663 -2587 1697 -2573
rect 1759 -2587 1793 -2573
rect 2483 -2471 2517 -2457
rect 2579 -2471 2613 -2457
rect 2483 -2491 2497 -2471
rect 2497 -2491 2517 -2471
rect 2579 -2491 2599 -2471
rect 2599 -2491 2613 -2471
rect 2483 -2573 2497 -2553
rect 2497 -2573 2517 -2553
rect 2579 -2573 2599 -2553
rect 2599 -2573 2613 -2553
rect 2483 -2587 2517 -2573
rect 2579 -2587 2613 -2573
rect 3303 -2471 3337 -2457
rect 3399 -2471 3433 -2457
rect 3303 -2491 3317 -2471
rect 3317 -2491 3337 -2471
rect 3399 -2491 3419 -2471
rect 3419 -2491 3433 -2471
rect 3303 -2573 3317 -2553
rect 3317 -2573 3337 -2553
rect 3399 -2573 3419 -2553
rect 3419 -2573 3433 -2553
rect 3303 -2587 3337 -2573
rect 3399 -2587 3433 -2573
rect 4123 -2471 4157 -2457
rect 4219 -2471 4253 -2457
rect 4123 -2491 4137 -2471
rect 4137 -2491 4157 -2471
rect 4219 -2491 4239 -2471
rect 4239 -2491 4253 -2471
rect 4123 -2573 4137 -2553
rect 4137 -2573 4157 -2553
rect 4219 -2573 4239 -2553
rect 4239 -2573 4253 -2553
rect 4123 -2587 4157 -2573
rect 4219 -2587 4253 -2573
rect 4943 -2471 4977 -2457
rect 5039 -2471 5073 -2457
rect 4943 -2491 4957 -2471
rect 4957 -2491 4977 -2471
rect 5039 -2491 5059 -2471
rect 5059 -2491 5073 -2471
rect 4943 -2573 4957 -2553
rect 4957 -2573 4977 -2553
rect 5039 -2573 5059 -2553
rect 5059 -2573 5073 -2553
rect 4943 -2587 4977 -2573
rect 5039 -2587 5073 -2573
rect 5763 -2471 5797 -2457
rect 5859 -2471 5893 -2457
rect 5763 -2491 5777 -2471
rect 5777 -2491 5797 -2471
rect 5859 -2491 5879 -2471
rect 5879 -2491 5893 -2471
rect 5763 -2573 5777 -2553
rect 5777 -2573 5797 -2553
rect 5859 -2573 5879 -2553
rect 5879 -2573 5893 -2553
rect 5763 -2587 5797 -2573
rect 5859 -2587 5893 -2573
rect 6583 -2471 6617 -2457
rect 6679 -2471 6713 -2457
rect 6583 -2491 6597 -2471
rect 6597 -2491 6617 -2471
rect 6679 -2491 6699 -2471
rect 6699 -2491 6713 -2471
rect 6583 -2573 6597 -2553
rect 6597 -2573 6617 -2553
rect 6679 -2573 6699 -2553
rect 6699 -2573 6713 -2553
rect 6583 -2587 6617 -2573
rect 6679 -2587 6713 -2573
rect -797 -3291 -763 -3277
rect -701 -3291 -667 -3277
rect -797 -3311 -783 -3291
rect -783 -3311 -763 -3291
rect -701 -3311 -681 -3291
rect -681 -3311 -667 -3291
rect -797 -3393 -783 -3373
rect -783 -3393 -763 -3373
rect -701 -3393 -681 -3373
rect -681 -3393 -667 -3373
rect -797 -3407 -763 -3393
rect -701 -3407 -667 -3393
rect 23 -3291 57 -3277
rect 119 -3291 153 -3277
rect 23 -3311 37 -3291
rect 37 -3311 57 -3291
rect 119 -3311 139 -3291
rect 139 -3311 153 -3291
rect 23 -3393 37 -3373
rect 37 -3393 57 -3373
rect 119 -3393 139 -3373
rect 139 -3393 153 -3373
rect 23 -3407 57 -3393
rect 119 -3407 153 -3393
rect 843 -3291 877 -3277
rect 939 -3291 973 -3277
rect 843 -3311 857 -3291
rect 857 -3311 877 -3291
rect 939 -3311 959 -3291
rect 959 -3311 973 -3291
rect 843 -3393 857 -3373
rect 857 -3393 877 -3373
rect 939 -3393 959 -3373
rect 959 -3393 973 -3373
rect 843 -3407 877 -3393
rect 939 -3407 973 -3393
rect 1663 -3291 1697 -3277
rect 1759 -3291 1793 -3277
rect 1663 -3311 1677 -3291
rect 1677 -3311 1697 -3291
rect 1759 -3311 1779 -3291
rect 1779 -3311 1793 -3291
rect 1663 -3393 1677 -3373
rect 1677 -3393 1697 -3373
rect 1759 -3393 1779 -3373
rect 1779 -3393 1793 -3373
rect 1663 -3407 1697 -3393
rect 1759 -3407 1793 -3393
rect 2483 -3291 2517 -3277
rect 2579 -3291 2613 -3277
rect 2483 -3311 2497 -3291
rect 2497 -3311 2517 -3291
rect 2579 -3311 2599 -3291
rect 2599 -3311 2613 -3291
rect 2483 -3393 2497 -3373
rect 2497 -3393 2517 -3373
rect 2579 -3393 2599 -3373
rect 2599 -3393 2613 -3373
rect 2483 -3407 2517 -3393
rect 2579 -3407 2613 -3393
rect 3303 -3291 3337 -3277
rect 3399 -3291 3433 -3277
rect 3303 -3311 3317 -3291
rect 3317 -3311 3337 -3291
rect 3399 -3311 3419 -3291
rect 3419 -3311 3433 -3291
rect 3303 -3393 3317 -3373
rect 3317 -3393 3337 -3373
rect 3399 -3393 3419 -3373
rect 3419 -3393 3433 -3373
rect 3303 -3407 3337 -3393
rect 3399 -3407 3433 -3393
rect 4123 -3291 4157 -3277
rect 4219 -3291 4253 -3277
rect 4123 -3311 4137 -3291
rect 4137 -3311 4157 -3291
rect 4219 -3311 4239 -3291
rect 4239 -3311 4253 -3291
rect 4123 -3393 4137 -3373
rect 4137 -3393 4157 -3373
rect 4219 -3393 4239 -3373
rect 4239 -3393 4253 -3373
rect 4123 -3407 4157 -3393
rect 4219 -3407 4253 -3393
rect 4943 -3291 4977 -3277
rect 5039 -3291 5073 -3277
rect 4943 -3311 4957 -3291
rect 4957 -3311 4977 -3291
rect 5039 -3311 5059 -3291
rect 5059 -3311 5073 -3291
rect 4943 -3393 4957 -3373
rect 4957 -3393 4977 -3373
rect 5039 -3393 5059 -3373
rect 5059 -3393 5073 -3373
rect 4943 -3407 4977 -3393
rect 5039 -3407 5073 -3393
rect 5763 -3291 5797 -3277
rect 5859 -3291 5893 -3277
rect 5763 -3311 5777 -3291
rect 5777 -3311 5797 -3291
rect 5859 -3311 5879 -3291
rect 5879 -3311 5893 -3291
rect 5763 -3393 5777 -3373
rect 5777 -3393 5797 -3373
rect 5859 -3393 5879 -3373
rect 5879 -3393 5893 -3373
rect 5763 -3407 5797 -3393
rect 5859 -3407 5893 -3393
rect 6583 -3291 6617 -3277
rect 6679 -3291 6713 -3277
rect 6583 -3311 6597 -3291
rect 6597 -3311 6617 -3291
rect 6679 -3311 6699 -3291
rect 6699 -3311 6713 -3291
rect 6583 -3393 6597 -3373
rect 6597 -3393 6617 -3373
rect 6679 -3393 6699 -3373
rect 6699 -3393 6713 -3373
rect 6583 -3407 6617 -3393
rect 6679 -3407 6713 -3393
rect -797 -4111 -763 -4097
rect -701 -4111 -667 -4097
rect -797 -4131 -783 -4111
rect -783 -4131 -763 -4111
rect -701 -4131 -681 -4111
rect -681 -4131 -667 -4111
rect -797 -4213 -783 -4193
rect -783 -4213 -763 -4193
rect -701 -4213 -681 -4193
rect -681 -4213 -667 -4193
rect -797 -4227 -763 -4213
rect -701 -4227 -667 -4213
rect 23 -4111 57 -4097
rect 119 -4111 153 -4097
rect 23 -4131 37 -4111
rect 37 -4131 57 -4111
rect 119 -4131 139 -4111
rect 139 -4131 153 -4111
rect 23 -4213 37 -4193
rect 37 -4213 57 -4193
rect 119 -4213 139 -4193
rect 139 -4213 153 -4193
rect 23 -4227 57 -4213
rect 119 -4227 153 -4213
rect 843 -4111 877 -4097
rect 939 -4111 973 -4097
rect 843 -4131 857 -4111
rect 857 -4131 877 -4111
rect 939 -4131 959 -4111
rect 959 -4131 973 -4111
rect 843 -4213 857 -4193
rect 857 -4213 877 -4193
rect 939 -4213 959 -4193
rect 959 -4213 973 -4193
rect 843 -4227 877 -4213
rect 939 -4227 973 -4213
rect 1663 -4111 1697 -4097
rect 1759 -4111 1793 -4097
rect 1663 -4131 1677 -4111
rect 1677 -4131 1697 -4111
rect 1759 -4131 1779 -4111
rect 1779 -4131 1793 -4111
rect 1663 -4213 1677 -4193
rect 1677 -4213 1697 -4193
rect 1759 -4213 1779 -4193
rect 1779 -4213 1793 -4193
rect 1663 -4227 1697 -4213
rect 1759 -4227 1793 -4213
rect 2483 -4111 2517 -4097
rect 2579 -4111 2613 -4097
rect 2483 -4131 2497 -4111
rect 2497 -4131 2517 -4111
rect 2579 -4131 2599 -4111
rect 2599 -4131 2613 -4111
rect 2483 -4213 2497 -4193
rect 2497 -4213 2517 -4193
rect 2579 -4213 2599 -4193
rect 2599 -4213 2613 -4193
rect 2483 -4227 2517 -4213
rect 2579 -4227 2613 -4213
rect 3303 -4111 3337 -4097
rect 3399 -4111 3433 -4097
rect 3303 -4131 3317 -4111
rect 3317 -4131 3337 -4111
rect 3399 -4131 3419 -4111
rect 3419 -4131 3433 -4111
rect 3303 -4213 3317 -4193
rect 3317 -4213 3337 -4193
rect 3399 -4213 3419 -4193
rect 3419 -4213 3433 -4193
rect 3303 -4227 3337 -4213
rect 3399 -4227 3433 -4213
rect 4123 -4111 4157 -4097
rect 4219 -4111 4253 -4097
rect 4123 -4131 4137 -4111
rect 4137 -4131 4157 -4111
rect 4219 -4131 4239 -4111
rect 4239 -4131 4253 -4111
rect 4123 -4213 4137 -4193
rect 4137 -4213 4157 -4193
rect 4219 -4213 4239 -4193
rect 4239 -4213 4253 -4193
rect 4123 -4227 4157 -4213
rect 4219 -4227 4253 -4213
rect 4943 -4111 4977 -4097
rect 5039 -4111 5073 -4097
rect 4943 -4131 4957 -4111
rect 4957 -4131 4977 -4111
rect 5039 -4131 5059 -4111
rect 5059 -4131 5073 -4111
rect 4943 -4213 4957 -4193
rect 4957 -4213 4977 -4193
rect 5039 -4213 5059 -4193
rect 5059 -4213 5073 -4193
rect 4943 -4227 4977 -4213
rect 5039 -4227 5073 -4213
rect 5763 -4111 5797 -4097
rect 5859 -4111 5893 -4097
rect 5763 -4131 5777 -4111
rect 5777 -4131 5797 -4111
rect 5859 -4131 5879 -4111
rect 5879 -4131 5893 -4111
rect 5763 -4213 5777 -4193
rect 5777 -4213 5797 -4193
rect 5859 -4213 5879 -4193
rect 5879 -4213 5893 -4193
rect 5763 -4227 5797 -4213
rect 5859 -4227 5893 -4213
rect 6583 -4111 6617 -4097
rect 6679 -4111 6713 -4097
rect 6583 -4131 6597 -4111
rect 6597 -4131 6617 -4111
rect 6679 -4131 6699 -4111
rect 6699 -4131 6713 -4111
rect 6583 -4213 6597 -4193
rect 6597 -4213 6617 -4193
rect 6679 -4213 6699 -4193
rect 6699 -4213 6713 -4193
rect 6583 -4227 6617 -4213
rect 6679 -4227 6713 -4213
<< metal1 >>
rect 7400 6240 7960 6270
rect 7400 5710 7560 6240
rect 6690 4800 7560 5710
rect 6690 4400 6780 4420
rect 6690 4360 6720 4400
rect 6760 4360 6780 4400
rect 6690 4340 6780 4360
rect 7400 4300 7560 4800
rect 7600 4300 7660 6240
rect 7700 4300 7760 6240
rect 7800 5710 7960 6240
rect 8320 6210 8790 6240
rect 8320 5710 8350 6210
rect 7800 4830 8350 5710
rect 8480 5680 9210 6210
rect 8490 5300 9210 5680
rect 8490 4830 8520 5300
rect 7800 4800 8520 4830
rect 8810 4840 9100 4920
rect 7800 4300 7960 4800
rect 8810 4710 8890 4840
rect 8050 4690 8890 4710
rect 8050 4650 8070 4690
rect 8110 4650 8890 4690
rect 8050 4630 8890 4650
rect 9080 4400 9340 4590
rect 15560 4400 16050 4590
rect 7400 4270 7960 4300
rect 7250 4190 7880 4210
rect 7250 4150 7500 4190
rect 7540 4150 7820 4190
rect 7860 4150 7880 4190
rect 7250 4130 7880 4150
rect 7250 4090 7330 4130
rect 6690 4010 7330 4090
rect 7400 4030 7960 4060
rect 6690 3960 7320 3980
rect 6690 3920 7260 3960
rect 7300 3920 7320 3960
rect 6690 3900 7320 3920
rect 6660 3520 6990 3550
rect 6660 2660 6860 3520
rect 6960 2660 6990 3520
rect 6660 2630 6990 2660
rect 7400 2570 7560 4030
rect 6540 2490 7560 2570
rect 7400 2090 7560 2490
rect 7600 2090 7660 4030
rect 7700 2090 7760 4030
rect 7800 2090 7960 4030
rect 8590 4040 9090 4070
rect 8590 3550 8620 4040
rect 8060 3520 8620 3550
rect 8060 2660 8100 3520
rect 8200 2660 8620 3520
rect 8760 3150 9090 4040
rect 20360 3800 22950 3880
rect 15590 3250 15740 3390
rect 8760 2660 8790 3150
rect 12080 2910 16150 2940
rect 12080 2830 12110 2910
rect 12490 2830 15740 2910
rect 16120 2830 16150 2910
rect 12080 2800 16150 2830
rect 17000 2910 17440 3580
rect 19610 3500 20050 3580
rect 17000 2830 17030 2910
rect 17410 2830 17440 2910
rect 17000 2800 17440 2830
rect 8060 2630 8790 2660
rect 7400 2060 7960 2090
rect 8320 2500 9090 2570
rect 15820 2560 16210 2570
rect 16240 2560 16250 2600
rect 8320 2470 9110 2500
rect 8320 1690 8350 2470
rect 8490 1690 9190 2470
rect 8320 1660 9190 1690
rect 15810 1660 16250 2560
rect 15820 1260 15940 1280
rect 15820 1220 15880 1260
rect 15920 1220 15940 1260
rect 15820 1200 15940 1220
rect 15990 1200 16250 1280
rect 15990 950 16070 1200
rect 9080 760 9340 950
rect 15560 930 16070 950
rect 15560 780 15850 930
rect 15920 780 16070 930
rect 15560 760 16070 780
rect 16210 760 16470 950
rect 22690 760 22950 950
rect 7240 610 7730 630
rect 7240 570 7260 610
rect 7300 570 7670 610
rect 7710 570 7730 610
rect 7240 550 7730 570
rect 6620 420 6760 450
rect 6620 40 6650 420
rect 6730 40 6760 420
rect 6620 -780 6760 40
rect -1110 -817 6760 -780
rect 7820 420 7960 450
rect 7820 40 7850 420
rect 7930 40 7960 420
rect 7820 -790 7960 40
rect 8590 380 9100 410
rect 8590 -480 8620 380
rect 8760 -480 9100 380
rect 8590 -510 9100 -480
rect 15780 -510 16220 410
rect -1110 -851 -797 -817
rect -763 -851 -701 -817
rect -667 -851 23 -817
rect 57 -851 119 -817
rect 153 -851 843 -817
rect 877 -851 939 -817
rect 973 -851 1663 -817
rect 1697 -851 1759 -817
rect 1793 -851 2483 -817
rect 2517 -851 2579 -817
rect 2613 -851 3303 -817
rect 3337 -851 3399 -817
rect 3433 -851 4123 -817
rect 4157 -851 4219 -817
rect 4253 -851 4943 -817
rect 4977 -851 5039 -817
rect 5073 -851 5763 -817
rect 5797 -851 5859 -817
rect 5893 -851 6583 -817
rect 6617 -851 6679 -817
rect 6713 -851 6760 -817
rect -1110 -913 6760 -851
rect -1110 -947 -797 -913
rect -763 -947 -701 -913
rect -667 -947 23 -913
rect 57 -947 119 -913
rect 153 -947 843 -913
rect 877 -947 939 -913
rect 973 -947 1663 -913
rect 1697 -947 1759 -913
rect 1793 -947 2483 -913
rect 2517 -947 2579 -913
rect 2613 -947 3303 -913
rect 3337 -947 3399 -913
rect 3433 -947 4123 -913
rect 4157 -947 4219 -913
rect 4253 -947 4943 -913
rect 4977 -947 5039 -913
rect 5073 -947 5763 -913
rect 5797 -947 5859 -913
rect 5893 -947 6583 -913
rect 6617 -947 6679 -913
rect 6713 -947 6760 -913
rect -1110 -1000 6760 -947
rect 7410 -817 7960 -790
rect 7410 -851 7433 -817
rect 7467 -851 7529 -817
rect 7563 -851 7960 -817
rect 7410 -913 7960 -851
rect 16130 -790 16210 -510
rect 16130 -870 17110 -790
rect 7410 -947 7433 -913
rect 7467 -947 7529 -913
rect 7563 -947 7960 -913
rect 7410 -970 7960 -947
rect 16970 -930 17110 -870
rect -1110 -1637 6740 -1000
rect -1110 -1671 -797 -1637
rect -763 -1671 -701 -1637
rect -667 -1671 23 -1637
rect 57 -1671 119 -1637
rect 153 -1671 843 -1637
rect 877 -1671 939 -1637
rect 973 -1671 1663 -1637
rect 1697 -1671 1759 -1637
rect 1793 -1671 2483 -1637
rect 2517 -1671 2579 -1637
rect 2613 -1671 3303 -1637
rect 3337 -1671 3399 -1637
rect 3433 -1671 4123 -1637
rect 4157 -1671 4219 -1637
rect 4253 -1671 4943 -1637
rect 4977 -1671 5039 -1637
rect 5073 -1671 5763 -1637
rect 5797 -1671 5859 -1637
rect 5893 -1671 6583 -1637
rect 6617 -1671 6679 -1637
rect 6713 -1671 6740 -1637
rect 8590 -1170 8790 -1140
rect 8590 -1630 8620 -1170
rect 8760 -1630 8790 -1170
rect 16970 -1310 17000 -930
rect 17080 -1310 17110 -930
rect 16970 -1340 17110 -1310
rect 8590 -1660 8790 -1630
rect -1110 -1733 6740 -1671
rect -1110 -1767 -797 -1733
rect -763 -1767 -701 -1733
rect -667 -1767 23 -1733
rect 57 -1767 119 -1733
rect 153 -1767 843 -1733
rect 877 -1767 939 -1733
rect 973 -1767 1663 -1733
rect 1697 -1767 1759 -1733
rect 1793 -1767 2483 -1733
rect 2517 -1767 2579 -1733
rect 2613 -1767 3303 -1733
rect 3337 -1767 3399 -1733
rect 3433 -1767 4123 -1733
rect 4157 -1767 4219 -1733
rect 4253 -1767 4943 -1733
rect 4977 -1767 5039 -1733
rect 5073 -1767 5763 -1733
rect 5797 -1767 5859 -1733
rect 5893 -1767 6583 -1733
rect 6617 -1767 6679 -1733
rect 6713 -1767 6740 -1733
rect -1110 -2457 6740 -1767
rect -1110 -2491 -797 -2457
rect -763 -2491 -701 -2457
rect -667 -2491 23 -2457
rect 57 -2491 119 -2457
rect 153 -2491 843 -2457
rect 877 -2491 939 -2457
rect 973 -2491 1663 -2457
rect 1697 -2491 1759 -2457
rect 1793 -2491 2483 -2457
rect 2517 -2491 2579 -2457
rect 2613 -2491 3303 -2457
rect 3337 -2491 3399 -2457
rect 3433 -2491 4123 -2457
rect 4157 -2491 4219 -2457
rect 4253 -2491 4943 -2457
rect 4977 -2491 5039 -2457
rect 5073 -2491 5763 -2457
rect 5797 -2491 5859 -2457
rect 5893 -2491 6583 -2457
rect 6617 -2491 6679 -2457
rect 6713 -2491 6740 -2457
rect -1110 -2553 6740 -2491
rect -1110 -2587 -797 -2553
rect -763 -2587 -701 -2553
rect -667 -2587 23 -2553
rect 57 -2587 119 -2553
rect 153 -2587 843 -2553
rect 877 -2587 939 -2553
rect 973 -2587 1663 -2553
rect 1697 -2587 1759 -2553
rect 1793 -2587 2483 -2553
rect 2517 -2587 2579 -2553
rect 2613 -2587 3303 -2553
rect 3337 -2587 3399 -2553
rect 3433 -2587 4123 -2553
rect 4157 -2587 4219 -2553
rect 4253 -2587 4943 -2553
rect 4977 -2587 5039 -2553
rect 5073 -2587 5763 -2553
rect 5797 -2587 5859 -2553
rect 5893 -2587 6583 -2553
rect 6617 -2587 6679 -2553
rect 6713 -2587 6740 -2553
rect -1110 -3277 6740 -2587
rect -1110 -3311 -797 -3277
rect -763 -3311 -701 -3277
rect -667 -3311 23 -3277
rect 57 -3311 119 -3277
rect 153 -3311 843 -3277
rect 877 -3311 939 -3277
rect 973 -3311 1663 -3277
rect 1697 -3311 1759 -3277
rect 1793 -3311 2483 -3277
rect 2517 -3311 2579 -3277
rect 2613 -3311 3303 -3277
rect 3337 -3311 3399 -3277
rect 3433 -3311 4123 -3277
rect 4157 -3311 4219 -3277
rect 4253 -3311 4943 -3277
rect 4977 -3311 5039 -3277
rect 5073 -3311 5763 -3277
rect 5797 -3311 5859 -3277
rect 5893 -3311 6583 -3277
rect 6617 -3311 6679 -3277
rect 6713 -3311 6740 -3277
rect -1110 -3373 6740 -3311
rect -1110 -3407 -797 -3373
rect -763 -3407 -701 -3373
rect -667 -3407 23 -3373
rect 57 -3407 119 -3373
rect 153 -3407 843 -3373
rect 877 -3407 939 -3373
rect 973 -3407 1663 -3373
rect 1697 -3407 1759 -3373
rect 1793 -3407 2483 -3373
rect 2517 -3407 2579 -3373
rect 2613 -3407 3303 -3373
rect 3337 -3407 3399 -3373
rect 3433 -3407 4123 -3373
rect 4157 -3407 4219 -3373
rect 4253 -3407 4943 -3373
rect 4977 -3407 5039 -3373
rect 5073 -3407 5763 -3373
rect 5797 -3407 5859 -3373
rect 5893 -3407 6583 -3373
rect 6617 -3407 6679 -3373
rect 6713 -3407 6740 -3373
rect -1110 -4097 6740 -3407
rect -1110 -4131 -797 -4097
rect -763 -4131 -701 -4097
rect -667 -4131 23 -4097
rect 57 -4131 119 -4097
rect 153 -4131 843 -4097
rect 877 -4131 939 -4097
rect 973 -4131 1663 -4097
rect 1697 -4131 1759 -4097
rect 1793 -4131 2483 -4097
rect 2517 -4131 2579 -4097
rect 2613 -4131 3303 -4097
rect 3337 -4131 3399 -4097
rect 3433 -4131 4123 -4097
rect 4157 -4131 4219 -4097
rect 4253 -4131 4943 -4097
rect 4977 -4131 5039 -4097
rect 5073 -4131 5763 -4097
rect 5797 -4131 5859 -4097
rect 5893 -4131 6583 -4097
rect 6617 -4131 6679 -4097
rect 6713 -4131 6740 -4097
rect -1110 -4193 6740 -4131
rect -1110 -4227 -797 -4193
rect -763 -4227 -701 -4193
rect -667 -4227 23 -4193
rect 57 -4227 119 -4193
rect 153 -4227 843 -4193
rect 877 -4227 939 -4193
rect 973 -4227 1663 -4193
rect 1697 -4227 1759 -4193
rect 1793 -4227 2483 -4193
rect 2517 -4227 2579 -4193
rect 2613 -4227 3303 -4193
rect 3337 -4227 3399 -4193
rect 3433 -4227 4123 -4193
rect 4157 -4227 4219 -4193
rect 4253 -4227 4943 -4193
rect 4977 -4227 5039 -4193
rect 5073 -4227 5763 -4193
rect 5797 -4227 5859 -4193
rect 5893 -4227 6583 -4193
rect 6617 -4227 6679 -4193
rect 6713 -4227 6740 -4193
rect -1110 -4260 6740 -4227
rect 8320 -3470 9040 -3440
rect 8320 -4320 8350 -3470
rect 8490 -4320 9040 -3470
rect 8320 -4350 9040 -4320
rect 9010 -5250 9270 -5060
rect 15490 -5250 15980 -5060
rect 8590 -5610 9020 -5580
rect 8590 -6470 8620 -5610
rect 8760 -6470 9020 -5610
rect 20320 -5850 22950 -5770
rect 8590 -6500 9020 -6470
<< via1 >>
rect 8350 5680 8480 6210
rect 8350 4830 8490 5680
rect 6860 2660 6960 3520
rect 8100 2660 8200 3520
rect 8620 2910 8760 4040
rect 8620 2830 8650 2910
rect 8650 2830 8730 2910
rect 8730 2830 8760 2910
rect 8620 2660 8760 2830
rect 8350 1690 8490 2470
rect 8620 -480 8760 380
rect 8620 -1630 8760 -1170
rect 8350 -4320 8490 -3470
rect 8620 -6470 8760 -5610
<< metal2 >>
rect 8320 6210 8520 6420
rect 8320 4830 8350 6210
rect 8480 5680 8520 6210
rect 8490 4830 8520 5680
rect 6830 3520 8230 3550
rect 6830 2660 6860 3520
rect 6960 2660 8100 3520
rect 8200 2660 8230 3520
rect 6830 2630 8230 2660
rect 8320 2470 8520 4830
rect 8320 1690 8350 2470
rect 8490 1690 8520 2470
rect 8320 -3470 8520 1690
rect 8320 -4320 8350 -3470
rect 8490 -4320 8520 -3470
rect 8320 -6640 8520 -4320
rect 8590 4040 8790 6420
rect 8590 2660 8620 4040
rect 8760 2660 8790 4040
rect 8590 380 8790 2660
rect 8590 -480 8620 380
rect 8760 -480 8790 380
rect 8590 -1170 8790 -480
rect 8590 -1630 8620 -1170
rect 8760 -1630 8790 -1170
rect 8590 -5610 8790 -1630
rect 8590 -6470 8620 -5610
rect 8760 -6470 8790 -5610
rect 8590 -6640 8790 -6470
use opamp  opamp_1
timestamp 1620822988
transform 1 0 9470 0 1 -6700
box -460 60 10850 3400
use opamp  opamp_0
timestamp 1620822988
transform 1 0 9540 0 1 2950
box -460 60 10850 3400
use opamp_square  opamp_square_0
timestamp 1620667237
transform 1 0 410 0 1 2450
box -460 -2450 6280 3400
use opamp_square  opamp_square_1
timestamp 1620667237
transform 1 0 9540 0 1 -690
box -460 -2450 6280 3400
use opamp_square  opamp_square_2
timestamp 1620667237
transform 1 0 16670 0 1 -690
box -460 -2450 6280 3400
<< labels >>
rlabel metal1 6840 3900 6970 3980 5 net4
rlabel metal1 6840 4010 6970 4090 5 net2
rlabel locali 6700 4200 6780 4300 3 net6
rlabel metal1 6620 -120 6760 -30 3 net1
rlabel metal2 8590 6350 8790 6420 1 gnd
rlabel metal2 8320 6350 8520 6420 1 vdd
rlabel metal1 8990 4840 9070 4920 1 net3
<< end >>
