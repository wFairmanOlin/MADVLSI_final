magic
tech sky130A
timestamp 1620787459
<< poly >>
rect 6280 1075 6320 1090
rect 6240 720 6280 730
rect 6240 700 6250 720
rect 6270 700 6280 720
rect 6240 690 6280 700
rect 5885 530 5890 545
rect 6275 480 6320 500
rect 5890 465 5895 480
rect 6240 250 6280 260
rect 6240 230 6250 250
rect 6270 230 6280 250
rect 6240 220 6280 230
<< polycont >>
rect 6250 700 6270 720
rect 6250 230 6270 250
<< locali >>
rect 5010 4730 6490 4750
rect 6430 1015 6450 4730
rect 6320 995 6450 1015
rect 6240 720 6280 730
rect 6240 700 6250 720
rect 6270 700 6295 720
rect 6240 690 6280 700
rect 6240 250 6280 260
rect 5870 225 5910 235
rect 5870 205 5880 225
rect 5900 205 5910 225
rect 6240 230 6250 250
rect 6270 240 6280 250
rect 6375 245 6415 255
rect 6375 240 6385 245
rect 6270 230 6300 240
rect 6240 220 6300 230
rect 6320 225 6385 240
rect 6405 225 6510 245
rect 6320 220 6415 225
rect 6375 215 6415 220
rect 5870 195 5910 205
rect 5890 50 5910 60
rect 5890 30 10610 50
<< viali >>
rect 5880 205 5900 225
rect 6385 225 6405 245
<< metal1 >>
rect 10585 4895 10590 4915
rect 6320 1575 6365 1580
rect 6320 1540 6325 1575
rect 6360 1540 6365 1575
rect 6320 1535 6365 1540
rect 6065 1180 6535 1270
rect 6375 245 6415 255
rect 5865 235 5915 240
rect 5865 195 5870 235
rect 5910 195 5915 235
rect 5865 190 5915 195
rect 6375 225 6385 245
rect 6405 225 6415 245
rect 6375 175 6415 225
rect 6370 170 6420 175
rect 6370 130 6375 170
rect 6415 130 6420 170
rect 6370 125 6420 130
rect 10580 130 10590 160
<< via1 >>
rect 6325 1540 6360 1575
rect 5870 225 5910 235
rect 5870 205 5880 225
rect 5880 205 5900 225
rect 5900 205 5910 225
rect 5870 195 5910 205
rect 6375 130 6415 170
rect 6600 125 6640 165
<< metal2 >>
rect 6320 1575 6415 1580
rect 6320 1540 6325 1575
rect 6360 1540 6415 1575
rect 6320 1535 6415 1540
rect 6370 435 6415 1535
rect 6370 430 6500 435
rect 6155 395 6500 430
rect 5865 235 5915 240
rect 5865 195 5870 235
rect 5910 195 5915 235
rect 5865 190 5915 195
rect 6370 170 6420 175
rect 6370 130 6375 170
rect 6415 130 6420 170
rect 6370 125 6420 130
rect 6460 165 6500 395
rect 6590 165 6645 170
rect 6460 125 6600 165
rect 6640 125 6645 165
rect 6590 120 6645 125
<< via2 >>
rect 6325 1540 6360 1575
rect 5870 195 5910 235
rect 6375 130 6415 170
<< metal3 >>
rect 6240 1575 6510 1580
rect 6285 1540 6325 1575
rect 6360 1540 6510 1575
rect 6285 1535 6510 1540
rect 5865 235 5915 240
rect 5865 195 5870 235
rect 5910 195 5915 235
rect 5865 190 5915 195
rect 6370 170 6420 175
rect 6370 130 6375 170
rect 6415 130 6420 170
rect 6370 125 6420 130
rect 6600 125 6640 165
<< via3 >>
rect 5870 195 5910 235
rect 6375 130 6415 170
<< mimcap >>
rect 6600 125 6640 165
<< metal4 >>
rect 6250 1430 6285 1465
rect 5565 1395 6285 1430
rect 5565 240 5600 1395
rect 5565 235 5915 240
rect 5565 195 5870 235
rect 5910 195 5915 235
rect 5565 190 5915 195
rect 6370 170 6420 175
rect 6370 130 6375 170
rect 6415 130 6420 170
rect 6370 125 6420 130
rect 6375 80 6410 125
rect 6375 45 6505 80
use xor  xor_0
timestamp 1620784958
transform 0 -1 6275 1 0 545
box -495 -45 760 675
use 4pf_cap  4pf_cap_0
timestamp 1620530160
transform 1 0 6730 0 1 845
box -245 -800 3785 4275
use time_delay_2  time_delay_2_0
timestamp 1620783427
transform 1 0 6520 0 1 4745
box -30 -4660 4090 230
use 500fF_cap  500fF_cap_0
timestamp 1620530576
transform 0 -1 6225 1 0 1455
box -15 -60 2015 1215
<< labels >>
rlabel locali 5010 4740 5010 4740 7 Vclk
port 1 w
rlabel locali 10610 40 10610 40 3 Vpulse
port 2 e
rlabel metal1 10590 145 10590 145 3 VN
port 3 e
rlabel metal1 10590 4905 10590 4905 3 VP
port 4 e
rlabel metal1 6320 1185 6320 1185 5 VP
rlabel poly 5890 530 5890 530 5 net3
rlabel poly 5895 465 5895 465 5 net2
rlabel locali 6295 220 6295 220 5 net1
rlabel locali 6430 225 6430 225 5 net1
<< end >>
