magic
tech sky130A
timestamp 1620667237
<< nwell >>
rect -120 1150 3030 1670
<< nmos >>
rect 0 390 60 540
rect 110 390 170 540
rect 220 390 280 540
rect 330 390 390 540
rect 440 390 500 540
rect 550 390 610 540
rect 660 390 720 540
rect 770 390 830 540
rect 880 390 940 540
rect 990 390 1050 540
rect 1100 390 1160 540
rect 1210 390 1270 540
rect 1320 390 1380 540
rect 1530 390 1590 540
rect 1640 390 1700 540
rect 1750 390 1810 540
rect 1860 390 1920 540
rect 1970 390 2030 540
rect 2080 390 2140 540
rect 2190 390 2250 540
rect 2300 390 2360 540
rect 2410 390 2470 540
rect 2520 390 2580 540
rect 2630 390 2690 540
rect 2740 390 2800 540
rect 2850 390 2910 540
rect 0 70 60 220
rect 110 70 170 220
rect 220 70 280 220
rect 330 70 390 220
rect 440 70 500 220
rect 550 70 610 220
rect 660 70 720 220
rect 770 70 830 220
rect 880 70 940 220
rect 990 70 1050 220
rect 1100 70 1160 220
rect 1210 70 1270 220
rect 1320 70 1380 220
rect 1530 70 1590 220
rect 1640 70 1700 220
rect 1750 70 1810 220
rect 1860 70 1920 220
rect 1970 70 2030 220
rect 2080 70 2140 220
rect 2190 70 2250 220
rect 2300 70 2360 220
rect 2410 70 2470 220
rect 2520 70 2580 220
rect 2630 70 2690 220
rect 2740 70 2800 220
rect 2850 70 2910 220
<< pmos >>
rect 0 1500 60 1650
rect 110 1500 170 1650
rect 220 1500 280 1650
rect 330 1500 390 1650
rect 440 1500 500 1650
rect 550 1500 610 1650
rect 660 1500 720 1650
rect 770 1500 830 1650
rect 880 1500 940 1650
rect 990 1500 1050 1650
rect 1100 1500 1160 1650
rect 1210 1500 1270 1650
rect 1320 1500 1380 1650
rect 1530 1500 1590 1650
rect 1640 1500 1700 1650
rect 1750 1500 1810 1650
rect 1860 1500 1920 1650
rect 1970 1500 2030 1650
rect 2080 1500 2140 1650
rect 2190 1500 2250 1650
rect 2300 1500 2360 1650
rect 2410 1500 2470 1650
rect 2520 1500 2580 1650
rect 2630 1500 2690 1650
rect 2740 1500 2800 1650
rect 2850 1500 2910 1650
rect 0 1170 60 1320
rect 110 1170 170 1320
rect 220 1170 280 1320
rect 330 1170 390 1320
rect 440 1170 500 1320
rect 550 1170 610 1320
rect 660 1170 720 1320
rect 770 1170 830 1320
rect 880 1170 940 1320
rect 990 1170 1050 1320
rect 1100 1170 1160 1320
rect 1210 1170 1270 1320
rect 1320 1170 1380 1320
rect 1530 1170 1590 1320
rect 1640 1170 1700 1320
rect 1750 1170 1810 1320
rect 1860 1170 1920 1320
rect 1970 1170 2030 1320
rect 2080 1170 2140 1320
rect 2190 1170 2250 1320
rect 2300 1170 2360 1320
rect 2410 1170 2470 1320
rect 2520 1170 2580 1320
rect 2630 1170 2690 1320
rect 2740 1170 2800 1320
rect 2850 1170 2910 1320
<< ndiff >>
rect -50 525 0 540
rect -50 405 -35 525
rect -15 405 0 525
rect -50 390 0 405
rect 60 525 110 540
rect 60 405 75 525
rect 95 405 110 525
rect 60 390 110 405
rect 170 525 220 540
rect 170 405 185 525
rect 205 405 220 525
rect 170 390 220 405
rect 280 525 330 540
rect 280 405 295 525
rect 315 405 330 525
rect 280 390 330 405
rect 390 525 440 540
rect 390 405 405 525
rect 425 405 440 525
rect 390 390 440 405
rect 500 525 550 540
rect 500 405 515 525
rect 535 405 550 525
rect 500 390 550 405
rect 610 525 660 540
rect 610 405 625 525
rect 645 405 660 525
rect 610 390 660 405
rect 720 525 770 540
rect 720 405 735 525
rect 755 405 770 525
rect 720 390 770 405
rect 830 390 880 540
rect 940 525 990 540
rect 940 405 955 525
rect 975 405 990 525
rect 940 390 990 405
rect 1050 525 1100 540
rect 1050 405 1065 525
rect 1085 405 1100 525
rect 1050 390 1100 405
rect 1160 525 1210 540
rect 1160 405 1175 525
rect 1195 405 1210 525
rect 1160 390 1210 405
rect 1270 525 1320 540
rect 1270 405 1285 525
rect 1305 405 1320 525
rect 1270 390 1320 405
rect 1380 525 1430 540
rect 1480 525 1530 540
rect 1380 405 1395 525
rect 1415 405 1430 525
rect 1480 405 1495 525
rect 1515 405 1530 525
rect 1380 390 1430 405
rect 1480 390 1530 405
rect 1590 525 1640 540
rect 1590 405 1605 525
rect 1625 405 1640 525
rect 1590 390 1640 405
rect 1700 525 1750 540
rect 1700 405 1715 525
rect 1735 405 1750 525
rect 1700 390 1750 405
rect 1810 525 1860 540
rect 1810 405 1825 525
rect 1845 405 1860 525
rect 1810 390 1860 405
rect 1920 525 1970 540
rect 1920 405 1935 525
rect 1955 405 1970 525
rect 1920 390 1970 405
rect 2030 390 2080 540
rect 2140 525 2190 540
rect 2140 405 2155 525
rect 2175 405 2190 525
rect 2140 390 2190 405
rect 2250 525 2300 540
rect 2250 405 2265 525
rect 2285 405 2300 525
rect 2250 390 2300 405
rect 2360 525 2410 540
rect 2360 405 2375 525
rect 2395 405 2410 525
rect 2360 390 2410 405
rect 2470 525 2520 540
rect 2470 405 2485 525
rect 2505 405 2520 525
rect 2470 390 2520 405
rect 2580 525 2630 540
rect 2580 405 2595 525
rect 2615 405 2630 525
rect 2580 390 2630 405
rect 2690 525 2740 540
rect 2690 405 2705 525
rect 2725 405 2740 525
rect 2690 390 2740 405
rect 2800 525 2850 540
rect 2800 405 2815 525
rect 2835 405 2850 525
rect 2800 390 2850 405
rect 2910 525 2960 540
rect 2910 405 2925 525
rect 2945 405 2960 525
rect 2910 390 2960 405
rect -50 205 0 220
rect -50 85 -35 205
rect -15 85 0 205
rect -50 70 0 85
rect 60 205 110 220
rect 60 85 75 205
rect 95 85 110 205
rect 60 70 110 85
rect 170 205 220 220
rect 170 85 185 205
rect 205 85 220 205
rect 170 70 220 85
rect 280 205 330 220
rect 280 85 295 205
rect 315 85 330 205
rect 280 70 330 85
rect 390 205 440 220
rect 390 85 405 205
rect 425 85 440 205
rect 390 70 440 85
rect 500 205 550 220
rect 500 85 515 205
rect 535 85 550 205
rect 500 70 550 85
rect 610 205 660 220
rect 610 85 625 205
rect 645 85 660 205
rect 610 70 660 85
rect 720 205 770 220
rect 720 85 735 205
rect 755 85 770 205
rect 720 70 770 85
rect 830 70 880 220
rect 940 205 990 220
rect 940 85 955 205
rect 975 85 990 205
rect 940 70 990 85
rect 1050 205 1100 220
rect 1050 85 1065 205
rect 1085 85 1100 205
rect 1050 70 1100 85
rect 1160 205 1210 220
rect 1160 85 1175 205
rect 1195 85 1210 205
rect 1160 70 1210 85
rect 1270 205 1320 220
rect 1270 85 1285 205
rect 1305 85 1320 205
rect 1270 70 1320 85
rect 1380 205 1430 220
rect 1480 205 1530 220
rect 1380 85 1395 205
rect 1415 85 1430 205
rect 1480 85 1495 205
rect 1515 85 1530 205
rect 1380 70 1430 85
rect 1480 70 1530 85
rect 1590 205 1640 220
rect 1590 85 1605 205
rect 1625 85 1640 205
rect 1590 70 1640 85
rect 1700 205 1750 220
rect 1700 85 1715 205
rect 1735 85 1750 205
rect 1700 70 1750 85
rect 1810 205 1860 220
rect 1810 85 1825 205
rect 1845 85 1860 205
rect 1810 70 1860 85
rect 1920 205 1970 220
rect 1920 85 1935 205
rect 1955 85 1970 205
rect 1920 70 1970 85
rect 2030 70 2080 220
rect 2140 205 2190 220
rect 2140 85 2155 205
rect 2175 85 2190 205
rect 2140 70 2190 85
rect 2250 205 2300 220
rect 2250 85 2265 205
rect 2285 85 2300 205
rect 2250 70 2300 85
rect 2360 205 2410 220
rect 2360 85 2375 205
rect 2395 85 2410 205
rect 2360 70 2410 85
rect 2470 205 2520 220
rect 2470 85 2485 205
rect 2505 85 2520 205
rect 2470 70 2520 85
rect 2580 205 2630 220
rect 2580 85 2595 205
rect 2615 85 2630 205
rect 2580 70 2630 85
rect 2690 205 2740 220
rect 2690 85 2705 205
rect 2725 85 2740 205
rect 2690 70 2740 85
rect 2800 205 2850 220
rect 2800 85 2815 205
rect 2835 85 2850 205
rect 2800 70 2850 85
rect 2910 205 2960 220
rect 2910 85 2925 205
rect 2945 85 2960 205
rect 2910 70 2960 85
<< pdiff >>
rect -50 1635 0 1650
rect -50 1515 -35 1635
rect -15 1515 0 1635
rect -50 1500 0 1515
rect 60 1635 110 1650
rect 60 1515 75 1635
rect 95 1515 110 1635
rect 60 1500 110 1515
rect 170 1635 220 1650
rect 170 1515 185 1635
rect 205 1515 220 1635
rect 170 1500 220 1515
rect 280 1635 330 1650
rect 280 1515 295 1635
rect 315 1515 330 1635
rect 280 1500 330 1515
rect 390 1635 440 1650
rect 390 1515 405 1635
rect 425 1515 440 1635
rect 390 1500 440 1515
rect 500 1635 550 1650
rect 500 1515 515 1635
rect 535 1515 550 1635
rect 500 1500 550 1515
rect 610 1635 660 1650
rect 610 1515 625 1635
rect 645 1515 660 1635
rect 610 1500 660 1515
rect 720 1635 770 1650
rect 720 1515 735 1635
rect 755 1515 770 1635
rect 720 1500 770 1515
rect 830 1500 880 1650
rect 940 1635 990 1650
rect 940 1515 955 1635
rect 975 1515 990 1635
rect 940 1500 990 1515
rect 1050 1635 1100 1650
rect 1050 1515 1065 1635
rect 1085 1515 1100 1635
rect 1050 1500 1100 1515
rect 1160 1635 1210 1650
rect 1160 1515 1175 1635
rect 1195 1515 1210 1635
rect 1160 1500 1210 1515
rect 1270 1635 1320 1650
rect 1270 1515 1285 1635
rect 1305 1515 1320 1635
rect 1270 1500 1320 1515
rect 1380 1635 1430 1650
rect 1480 1635 1530 1650
rect 1380 1515 1395 1635
rect 1415 1515 1430 1635
rect 1480 1515 1495 1635
rect 1515 1515 1530 1635
rect 1380 1500 1430 1515
rect 1480 1500 1530 1515
rect 1590 1635 1640 1650
rect 1590 1515 1605 1635
rect 1625 1515 1640 1635
rect 1590 1500 1640 1515
rect 1700 1635 1750 1650
rect 1700 1515 1715 1635
rect 1735 1515 1750 1635
rect 1700 1500 1750 1515
rect 1810 1635 1860 1650
rect 1810 1515 1825 1635
rect 1845 1515 1860 1635
rect 1810 1500 1860 1515
rect 1920 1635 1970 1650
rect 1920 1515 1935 1635
rect 1955 1515 1970 1635
rect 1920 1500 1970 1515
rect 2030 1500 2080 1650
rect 2140 1635 2190 1650
rect 2140 1515 2155 1635
rect 2175 1515 2190 1635
rect 2140 1500 2190 1515
rect 2250 1635 2300 1650
rect 2250 1515 2265 1635
rect 2285 1515 2300 1635
rect 2250 1500 2300 1515
rect 2360 1635 2410 1650
rect 2360 1515 2375 1635
rect 2395 1515 2410 1635
rect 2360 1500 2410 1515
rect 2470 1635 2520 1650
rect 2470 1515 2485 1635
rect 2505 1515 2520 1635
rect 2470 1500 2520 1515
rect 2580 1635 2630 1650
rect 2580 1515 2595 1635
rect 2615 1515 2630 1635
rect 2580 1500 2630 1515
rect 2690 1635 2740 1650
rect 2690 1515 2705 1635
rect 2725 1515 2740 1635
rect 2690 1500 2740 1515
rect 2800 1635 2850 1650
rect 2800 1515 2815 1635
rect 2835 1515 2850 1635
rect 2800 1500 2850 1515
rect 2910 1635 2960 1650
rect 2910 1515 2925 1635
rect 2945 1515 2960 1635
rect 2910 1500 2960 1515
rect -50 1305 0 1320
rect -50 1185 -35 1305
rect -15 1185 0 1305
rect -50 1170 0 1185
rect 60 1305 110 1320
rect 60 1185 75 1305
rect 95 1185 110 1305
rect 60 1170 110 1185
rect 170 1305 220 1320
rect 170 1185 185 1305
rect 205 1185 220 1305
rect 170 1170 220 1185
rect 280 1305 330 1320
rect 280 1185 295 1305
rect 315 1185 330 1305
rect 280 1170 330 1185
rect 390 1305 440 1320
rect 390 1185 405 1305
rect 425 1185 440 1305
rect 390 1170 440 1185
rect 500 1305 550 1320
rect 500 1185 515 1305
rect 535 1185 550 1305
rect 500 1170 550 1185
rect 610 1305 660 1320
rect 610 1185 625 1305
rect 645 1185 660 1305
rect 610 1170 660 1185
rect 720 1305 770 1320
rect 720 1185 735 1305
rect 755 1185 770 1305
rect 720 1170 770 1185
rect 830 1170 880 1320
rect 940 1305 990 1320
rect 940 1185 955 1305
rect 975 1185 990 1305
rect 940 1170 990 1185
rect 1050 1305 1100 1320
rect 1050 1185 1065 1305
rect 1085 1185 1100 1305
rect 1050 1170 1100 1185
rect 1160 1305 1210 1320
rect 1160 1185 1175 1305
rect 1195 1185 1210 1305
rect 1160 1170 1210 1185
rect 1270 1305 1320 1320
rect 1270 1185 1285 1305
rect 1305 1185 1320 1305
rect 1270 1170 1320 1185
rect 1380 1305 1430 1320
rect 1480 1305 1530 1320
rect 1380 1185 1395 1305
rect 1415 1185 1430 1305
rect 1480 1185 1495 1305
rect 1515 1185 1530 1305
rect 1380 1170 1430 1185
rect 1480 1170 1530 1185
rect 1590 1305 1640 1320
rect 1590 1185 1605 1305
rect 1625 1185 1640 1305
rect 1590 1170 1640 1185
rect 1700 1305 1750 1320
rect 1700 1185 1715 1305
rect 1735 1185 1750 1305
rect 1700 1170 1750 1185
rect 1810 1305 1860 1320
rect 1810 1185 1825 1305
rect 1845 1185 1860 1305
rect 1810 1170 1860 1185
rect 1920 1305 1970 1320
rect 1920 1185 1935 1305
rect 1955 1185 1970 1305
rect 1920 1170 1970 1185
rect 2030 1170 2080 1320
rect 2140 1305 2190 1320
rect 2140 1185 2155 1305
rect 2175 1185 2190 1305
rect 2140 1170 2190 1185
rect 2250 1305 2300 1320
rect 2250 1185 2265 1305
rect 2285 1185 2300 1305
rect 2250 1170 2300 1185
rect 2360 1305 2410 1320
rect 2360 1185 2375 1305
rect 2395 1185 2410 1305
rect 2360 1170 2410 1185
rect 2470 1305 2520 1320
rect 2470 1185 2485 1305
rect 2505 1185 2520 1305
rect 2470 1170 2520 1185
rect 2580 1305 2630 1320
rect 2580 1185 2595 1305
rect 2615 1185 2630 1305
rect 2580 1170 2630 1185
rect 2690 1305 2740 1320
rect 2690 1185 2705 1305
rect 2725 1185 2740 1305
rect 2690 1170 2740 1185
rect 2800 1305 2850 1320
rect 2800 1185 2815 1305
rect 2835 1185 2850 1305
rect 2800 1170 2850 1185
rect 2910 1305 2960 1320
rect 2910 1185 2925 1305
rect 2945 1185 2960 1305
rect 2910 1170 2960 1185
<< ndiffc >>
rect -35 405 -15 525
rect 75 405 95 525
rect 185 405 205 525
rect 295 405 315 525
rect 405 405 425 525
rect 515 405 535 525
rect 625 405 645 525
rect 735 405 755 525
rect 955 405 975 525
rect 1065 405 1085 525
rect 1175 405 1195 525
rect 1285 405 1305 525
rect 1395 405 1415 525
rect 1495 405 1515 525
rect 1605 405 1625 525
rect 1715 405 1735 525
rect 1825 405 1845 525
rect 1935 405 1955 525
rect 2155 405 2175 525
rect 2265 405 2285 525
rect 2375 405 2395 525
rect 2485 405 2505 525
rect 2595 405 2615 525
rect 2705 405 2725 525
rect 2815 405 2835 525
rect 2925 405 2945 525
rect -35 85 -15 205
rect 75 85 95 205
rect 185 85 205 205
rect 295 85 315 205
rect 405 85 425 205
rect 515 85 535 205
rect 625 85 645 205
rect 735 85 755 205
rect 955 85 975 205
rect 1065 85 1085 205
rect 1175 85 1195 205
rect 1285 85 1305 205
rect 1395 85 1415 205
rect 1495 85 1515 205
rect 1605 85 1625 205
rect 1715 85 1735 205
rect 1825 85 1845 205
rect 1935 85 1955 205
rect 2155 85 2175 205
rect 2265 85 2285 205
rect 2375 85 2395 205
rect 2485 85 2505 205
rect 2595 85 2615 205
rect 2705 85 2725 205
rect 2815 85 2835 205
rect 2925 85 2945 205
<< pdiffc >>
rect -35 1515 -15 1635
rect 75 1515 95 1635
rect 185 1515 205 1635
rect 295 1515 315 1635
rect 405 1515 425 1635
rect 515 1515 535 1635
rect 625 1515 645 1635
rect 735 1515 755 1635
rect 955 1515 975 1635
rect 1065 1515 1085 1635
rect 1175 1515 1195 1635
rect 1285 1515 1305 1635
rect 1395 1515 1415 1635
rect 1495 1515 1515 1635
rect 1605 1515 1625 1635
rect 1715 1515 1735 1635
rect 1825 1515 1845 1635
rect 1935 1515 1955 1635
rect 2155 1515 2175 1635
rect 2265 1515 2285 1635
rect 2375 1515 2395 1635
rect 2485 1515 2505 1635
rect 2595 1515 2615 1635
rect 2705 1515 2725 1635
rect 2815 1515 2835 1635
rect 2925 1515 2945 1635
rect -35 1185 -15 1305
rect 75 1185 95 1305
rect 185 1185 205 1305
rect 295 1185 315 1305
rect 405 1185 425 1305
rect 515 1185 535 1305
rect 625 1185 645 1305
rect 735 1185 755 1305
rect 955 1185 975 1305
rect 1065 1185 1085 1305
rect 1175 1185 1195 1305
rect 1285 1185 1305 1305
rect 1395 1185 1415 1305
rect 1495 1185 1515 1305
rect 1605 1185 1625 1305
rect 1715 1185 1735 1305
rect 1825 1185 1845 1305
rect 1935 1185 1955 1305
rect 2155 1185 2175 1305
rect 2265 1185 2285 1305
rect 2375 1185 2395 1305
rect 2485 1185 2505 1305
rect 2595 1185 2615 1305
rect 2705 1185 2725 1305
rect 2815 1185 2835 1305
rect 2925 1185 2945 1305
<< psubdiff >>
rect -100 525 -50 540
rect -100 405 -85 525
rect -65 405 -50 525
rect -100 390 -50 405
rect 1430 525 1480 540
rect 1430 405 1445 525
rect 1465 405 1480 525
rect 1430 390 1480 405
rect 2960 525 3010 540
rect 2960 405 2975 525
rect 2995 405 3010 525
rect 2960 390 3010 405
rect -100 205 -50 220
rect -100 85 -85 205
rect -65 85 -50 205
rect -100 70 -50 85
rect 1430 205 1480 220
rect 1430 85 1445 205
rect 1465 85 1480 205
rect 1430 70 1480 85
rect 2960 205 3010 220
rect 2960 85 2975 205
rect 2995 85 3010 205
rect 2960 70 3010 85
<< nsubdiff >>
rect -100 1635 -50 1650
rect -100 1515 -85 1635
rect -65 1515 -50 1635
rect -100 1500 -50 1515
rect 1430 1635 1480 1650
rect 1430 1515 1445 1635
rect 1465 1515 1480 1635
rect 1430 1500 1480 1515
rect 2960 1635 3010 1650
rect 2960 1515 2975 1635
rect 2995 1515 3010 1635
rect 2960 1500 3010 1515
rect -100 1305 -50 1320
rect -100 1185 -85 1305
rect -65 1185 -50 1305
rect -100 1170 -50 1185
rect 1430 1305 1480 1320
rect 1430 1185 1445 1305
rect 1465 1185 1480 1305
rect 1430 1170 1480 1185
rect 2960 1305 3010 1320
rect 2960 1185 2975 1305
rect 2995 1185 3010 1305
rect 2960 1170 3010 1185
<< psubdiffcont >>
rect -85 405 -65 525
rect 1445 405 1465 525
rect 2975 405 2995 525
rect -85 85 -65 205
rect 1445 85 1465 205
rect 2975 85 2995 205
<< nsubdiffcont >>
rect -85 1515 -65 1635
rect 1445 1515 1465 1635
rect 2975 1515 2995 1635
rect -85 1185 -65 1305
rect 1445 1185 1465 1305
rect 2975 1185 2995 1305
<< poly >>
rect 0 1650 60 1665
rect 110 1650 170 1665
rect 220 1650 280 1665
rect 330 1650 390 1665
rect 440 1650 500 1665
rect 550 1650 610 1665
rect 660 1650 720 1665
rect 770 1650 830 1665
rect 880 1650 940 1665
rect 990 1650 1050 1665
rect 1100 1650 1160 1665
rect 1210 1650 1270 1665
rect 1320 1650 1380 1665
rect 1530 1650 1590 1665
rect 1640 1650 1700 1665
rect 1750 1650 1810 1665
rect 1860 1650 1920 1665
rect 1970 1650 2030 1665
rect 2080 1650 2140 1665
rect 2190 1650 2250 1665
rect 2300 1650 2360 1665
rect 2410 1650 2470 1665
rect 2520 1650 2580 1665
rect 2630 1650 2690 1665
rect 2740 1650 2800 1665
rect 2850 1650 2910 1665
rect 0 1475 60 1500
rect 0 1455 20 1475
rect 40 1455 60 1475
rect 0 1320 60 1455
rect 110 1420 170 1500
rect 110 1400 130 1420
rect 150 1400 170 1420
rect 110 1320 170 1400
rect 220 1420 280 1500
rect 220 1400 240 1420
rect 260 1400 280 1420
rect 220 1390 280 1400
rect 330 1420 390 1500
rect 440 1485 500 1500
rect 550 1485 610 1500
rect 440 1475 610 1485
rect 440 1455 515 1475
rect 535 1455 610 1475
rect 440 1445 610 1455
rect 660 1475 720 1500
rect 660 1455 680 1475
rect 700 1455 720 1475
rect 660 1440 720 1455
rect 770 1485 830 1500
rect 880 1485 940 1500
rect 770 1475 940 1485
rect 770 1455 900 1475
rect 920 1455 940 1475
rect 770 1440 940 1455
rect 330 1400 350 1420
rect 370 1400 390 1420
rect 220 1320 280 1335
rect 330 1320 390 1400
rect 440 1365 500 1375
rect 440 1345 460 1365
rect 480 1345 500 1365
rect 440 1320 500 1345
rect 550 1365 610 1375
rect 550 1345 570 1365
rect 590 1345 610 1365
rect 550 1320 610 1345
rect 660 1320 720 1335
rect 770 1320 830 1440
rect 880 1320 940 1440
rect 990 1320 1050 1500
rect 1100 1420 1160 1500
rect 1100 1400 1120 1420
rect 1140 1400 1160 1420
rect 1100 1320 1160 1400
rect 1210 1320 1270 1500
rect 1320 1320 1380 1500
rect 1530 1320 1590 1500
rect 1640 1320 1700 1500
rect 1750 1420 1810 1500
rect 1750 1400 1770 1420
rect 1790 1400 1810 1420
rect 1750 1320 1810 1400
rect 1860 1320 1920 1500
rect 1970 1485 2030 1500
rect 2080 1485 2140 1500
rect 1970 1475 2140 1485
rect 1970 1455 1990 1475
rect 2010 1455 2140 1475
rect 1970 1440 2140 1455
rect 2190 1475 2250 1500
rect 2190 1455 2210 1475
rect 2230 1455 2250 1475
rect 2190 1440 2250 1455
rect 2300 1485 2360 1500
rect 2410 1485 2470 1500
rect 2300 1475 2470 1485
rect 2300 1455 2375 1475
rect 2395 1455 2470 1475
rect 2300 1445 2470 1455
rect 1970 1320 2030 1440
rect 2080 1320 2140 1440
rect 2520 1420 2580 1500
rect 2520 1400 2540 1420
rect 2560 1400 2580 1420
rect 2300 1365 2360 1375
rect 2300 1345 2320 1365
rect 2340 1345 2360 1365
rect 2190 1320 2250 1335
rect 2300 1320 2360 1345
rect 2410 1365 2470 1375
rect 2410 1345 2430 1365
rect 2450 1345 2470 1365
rect 2410 1320 2470 1345
rect 2520 1320 2580 1400
rect 2630 1420 2690 1500
rect 2630 1400 2650 1420
rect 2670 1400 2690 1420
rect 2630 1390 2690 1400
rect 2740 1420 2800 1500
rect 2740 1400 2760 1420
rect 2780 1400 2800 1420
rect 2630 1320 2690 1335
rect 2740 1320 2800 1400
rect 2850 1475 2910 1500
rect 2850 1455 2870 1475
rect 2890 1455 2910 1475
rect 2850 1320 2910 1455
rect 0 1150 60 1170
rect 110 1150 170 1170
rect 220 1145 280 1170
rect 330 1155 390 1170
rect 440 1155 500 1170
rect 550 1155 610 1170
rect 220 1125 240 1145
rect 260 1125 280 1145
rect 220 1110 280 1125
rect 660 1145 720 1170
rect 770 1150 830 1170
rect 880 1150 940 1170
rect 660 1125 680 1145
rect 700 1125 720 1145
rect 660 1110 720 1125
rect 990 1145 1050 1170
rect 1100 1150 1160 1170
rect 990 1125 1010 1145
rect 1030 1125 1050 1145
rect 990 1110 1050 1125
rect 1210 1145 1270 1170
rect 1210 1125 1230 1145
rect 1250 1125 1270 1145
rect 1210 1110 1270 1125
rect 1320 1145 1380 1170
rect 1320 1125 1340 1145
rect 1360 1125 1380 1145
rect 1320 1110 1380 1125
rect 1530 1145 1590 1170
rect 1530 1125 1550 1145
rect 1570 1125 1590 1145
rect 1530 1110 1590 1125
rect 1640 1145 1700 1170
rect 1750 1150 1810 1170
rect 1640 1125 1660 1145
rect 1680 1125 1700 1145
rect 1640 1110 1700 1125
rect 1860 1145 1920 1170
rect 1970 1150 2030 1170
rect 2080 1150 2140 1170
rect 1860 1125 1880 1145
rect 1900 1125 1920 1145
rect 1860 1110 1920 1125
rect 2190 1145 2250 1170
rect 2300 1155 2360 1170
rect 2410 1155 2470 1170
rect 2520 1155 2580 1170
rect 2190 1125 2210 1145
rect 2230 1125 2250 1145
rect 2190 1110 2250 1125
rect 2630 1145 2690 1170
rect 2740 1150 2800 1170
rect 2850 1150 2910 1170
rect 2630 1125 2650 1145
rect 2670 1125 2690 1145
rect 2630 1110 2690 1125
rect 220 580 280 595
rect 220 560 240 580
rect 260 560 280 580
rect 0 540 60 555
rect 110 540 170 555
rect 220 540 280 560
rect 660 580 720 595
rect 660 560 680 580
rect 700 560 720 580
rect 330 540 390 555
rect 440 540 500 555
rect 550 540 610 555
rect 660 540 720 560
rect 990 580 1050 595
rect 990 560 1010 580
rect 1030 560 1050 580
rect 770 540 830 555
rect 880 540 940 555
rect 990 540 1050 560
rect 1210 580 1270 595
rect 1210 560 1230 580
rect 1250 560 1270 580
rect 1100 540 1160 555
rect 1210 540 1270 560
rect 1320 580 1380 595
rect 1320 560 1340 580
rect 1360 560 1380 580
rect 1320 540 1380 560
rect 1530 580 1590 595
rect 1530 560 1550 580
rect 1570 560 1590 580
rect 1530 540 1590 560
rect 1640 580 1700 595
rect 1640 560 1660 580
rect 1680 560 1700 580
rect 1640 540 1700 560
rect 1860 580 1920 595
rect 1860 560 1880 580
rect 1900 560 1920 580
rect 1750 540 1810 555
rect 1860 540 1920 560
rect 2190 580 2250 595
rect 2190 560 2210 580
rect 2230 560 2250 580
rect 1970 540 2030 555
rect 2080 540 2140 555
rect 2190 540 2250 560
rect 2630 580 2690 595
rect 2630 560 2650 580
rect 2670 560 2690 580
rect 2300 540 2360 555
rect 2410 540 2470 555
rect 2520 540 2580 555
rect 2630 540 2690 560
rect 2740 540 2800 555
rect 2850 540 2910 555
rect 0 260 60 390
rect 0 240 20 260
rect 40 240 60 260
rect 0 220 60 240
rect 110 315 170 390
rect 220 375 280 390
rect 110 295 130 315
rect 150 295 170 315
rect 110 220 170 295
rect 220 315 280 325
rect 220 295 240 315
rect 260 295 280 315
rect 220 220 280 295
rect 330 315 390 390
rect 440 370 500 390
rect 440 350 460 370
rect 480 350 500 370
rect 440 340 500 350
rect 550 370 610 390
rect 660 375 720 390
rect 550 350 570 370
rect 590 350 610 370
rect 550 340 610 350
rect 330 295 350 315
rect 370 295 390 315
rect 330 220 390 295
rect 770 275 830 390
rect 880 275 940 390
rect 440 260 610 270
rect 440 240 515 260
rect 535 240 610 260
rect 440 230 610 240
rect 440 220 500 230
rect 550 220 610 230
rect 660 260 720 275
rect 660 240 680 260
rect 700 240 720 260
rect 660 220 720 240
rect 770 260 940 275
rect 770 240 900 260
rect 920 240 940 260
rect 770 230 940 240
rect 770 220 830 230
rect 880 220 940 230
rect 990 220 1050 390
rect 1100 315 1160 390
rect 1210 375 1270 390
rect 1100 295 1120 315
rect 1140 295 1160 315
rect 1100 220 1160 295
rect 1210 260 1270 275
rect 1210 240 1230 260
rect 1250 240 1270 260
rect 1210 220 1270 240
rect 1320 220 1380 390
rect 1530 220 1590 390
rect 1640 375 1700 390
rect 1750 315 1810 390
rect 1750 295 1770 315
rect 1790 295 1810 315
rect 1640 260 1700 275
rect 1640 240 1660 260
rect 1680 240 1700 260
rect 1640 220 1700 240
rect 1750 220 1810 295
rect 1860 220 1920 390
rect 1970 275 2030 390
rect 2080 275 2140 390
rect 2190 375 2250 390
rect 2300 370 2360 390
rect 2300 350 2320 370
rect 2340 350 2360 370
rect 2300 340 2360 350
rect 2410 370 2470 390
rect 2410 350 2430 370
rect 2450 350 2470 370
rect 2410 340 2470 350
rect 2520 315 2580 390
rect 2630 375 2690 390
rect 2520 295 2540 315
rect 2560 295 2580 315
rect 1970 260 2140 275
rect 1970 240 1990 260
rect 2010 240 2140 260
rect 1970 230 2140 240
rect 1970 220 2030 230
rect 2080 220 2140 230
rect 2190 260 2250 275
rect 2190 240 2210 260
rect 2230 240 2250 260
rect 2190 220 2250 240
rect 2300 260 2470 270
rect 2300 240 2375 260
rect 2395 240 2470 260
rect 2300 230 2470 240
rect 2300 220 2360 230
rect 2410 220 2470 230
rect 2520 220 2580 295
rect 2630 315 2690 325
rect 2630 295 2650 315
rect 2670 295 2690 315
rect 2630 220 2690 295
rect 2740 315 2800 390
rect 2740 295 2760 315
rect 2780 295 2800 315
rect 2740 220 2800 295
rect 2850 260 2910 390
rect 2850 240 2870 260
rect 2890 240 2910 260
rect 2850 220 2910 240
rect 0 55 60 70
rect 110 55 170 70
rect 220 55 280 70
rect 330 55 390 70
rect 440 55 500 70
rect 550 55 610 70
rect 660 55 720 70
rect 770 55 830 70
rect 880 55 940 70
rect 990 55 1050 70
rect 1100 55 1160 70
rect 1210 55 1270 70
rect 1320 55 1380 70
rect 1530 55 1590 70
rect 1640 55 1700 70
rect 1750 55 1810 70
rect 1860 55 1920 70
rect 1970 55 2030 70
rect 2080 55 2140 70
rect 2190 55 2250 70
rect 2300 55 2360 70
rect 2410 55 2470 70
rect 2520 55 2580 70
rect 2630 55 2690 70
rect 2740 55 2800 70
rect 2850 55 2910 70
<< polycont >>
rect 20 1455 40 1475
rect 130 1400 150 1420
rect 240 1400 260 1420
rect 515 1455 535 1475
rect 680 1455 700 1475
rect 900 1455 920 1475
rect 350 1400 370 1420
rect 460 1345 480 1365
rect 570 1345 590 1365
rect 1120 1400 1140 1420
rect 1770 1400 1790 1420
rect 1990 1455 2010 1475
rect 2210 1455 2230 1475
rect 2375 1455 2395 1475
rect 2540 1400 2560 1420
rect 2320 1345 2340 1365
rect 2430 1345 2450 1365
rect 2650 1400 2670 1420
rect 2760 1400 2780 1420
rect 2870 1455 2890 1475
rect 240 1125 260 1145
rect 680 1125 700 1145
rect 1010 1125 1030 1145
rect 1230 1125 1250 1145
rect 1340 1125 1360 1145
rect 1550 1125 1570 1145
rect 1660 1125 1680 1145
rect 1880 1125 1900 1145
rect 2210 1125 2230 1145
rect 2650 1125 2670 1145
rect 240 560 260 580
rect 680 560 700 580
rect 1010 560 1030 580
rect 1230 560 1250 580
rect 1340 560 1360 580
rect 1550 560 1570 580
rect 1660 560 1680 580
rect 1880 560 1900 580
rect 2210 560 2230 580
rect 2650 560 2670 580
rect 20 240 40 260
rect 130 295 150 315
rect 240 295 260 315
rect 460 350 480 370
rect 570 350 590 370
rect 350 295 370 315
rect 515 240 535 260
rect 680 240 700 260
rect 900 240 920 260
rect 1120 295 1140 315
rect 1230 240 1250 260
rect 1770 295 1790 315
rect 1660 240 1680 260
rect 2320 350 2340 370
rect 2430 350 2450 370
rect 2540 295 2560 315
rect 1990 240 2010 260
rect 2210 240 2230 260
rect 2375 240 2395 260
rect 2650 295 2670 315
rect 2760 295 2780 315
rect 2870 240 2890 260
<< locali >>
rect -215 1690 -175 1700
rect -215 1670 -205 1690
rect -185 1670 -175 1690
rect -215 525 -175 1670
rect 65 1690 105 1700
rect 65 1670 75 1690
rect 95 1670 105 1690
rect -95 1635 -5 1645
rect -95 1515 -85 1635
rect -65 1515 -35 1635
rect -15 1515 -5 1635
rect -95 1485 -5 1515
rect 65 1635 105 1670
rect 285 1690 325 1700
rect 285 1670 295 1690
rect 315 1670 325 1690
rect 65 1515 75 1635
rect 95 1515 105 1635
rect 65 1505 105 1515
rect 175 1635 215 1645
rect 175 1515 185 1635
rect 205 1515 215 1635
rect -95 1475 50 1485
rect -95 1455 20 1475
rect 40 1455 50 1475
rect -95 1445 50 1455
rect 175 1480 215 1515
rect 285 1635 325 1670
rect 2585 1690 2625 1700
rect 2585 1670 2595 1690
rect 2615 1670 2625 1690
rect 285 1515 295 1635
rect 315 1515 325 1635
rect 285 1505 325 1515
rect 395 1635 435 1645
rect 395 1515 405 1635
rect 425 1515 435 1635
rect 395 1505 435 1515
rect 505 1635 545 1645
rect 505 1515 515 1635
rect 535 1515 545 1635
rect 395 1480 430 1505
rect 175 1450 430 1480
rect -95 1305 -5 1445
rect 120 1420 270 1430
rect 120 1400 130 1420
rect 150 1400 185 1420
rect 205 1400 240 1420
rect 260 1400 270 1420
rect 120 1390 270 1400
rect 340 1420 380 1430
rect 340 1400 350 1420
rect 370 1400 380 1420
rect 340 1390 380 1400
rect -215 505 -205 525
rect -185 505 -175 525
rect -215 495 -175 505
rect -155 1205 -115 1215
rect -155 1185 -145 1205
rect -125 1185 -115 1205
rect -155 50 -115 1185
rect -95 1185 -85 1305
rect -65 1185 -35 1305
rect -15 1185 -5 1305
rect -95 1175 -5 1185
rect 65 1305 105 1315
rect 65 1185 75 1305
rect 95 1185 105 1305
rect 65 1175 105 1185
rect 175 1305 215 1390
rect 400 1315 430 1450
rect 505 1475 545 1515
rect 615 1635 655 1645
rect 615 1515 625 1635
rect 645 1515 655 1635
rect 615 1505 655 1515
rect 725 1635 765 1645
rect 725 1515 735 1635
rect 755 1535 765 1635
rect 945 1635 985 1645
rect 755 1515 870 1535
rect 725 1505 870 1515
rect 945 1515 955 1635
rect 975 1515 985 1635
rect 945 1505 985 1515
rect 1055 1635 1095 1645
rect 1055 1515 1065 1635
rect 1085 1515 1095 1635
rect 1055 1505 1095 1515
rect 1165 1635 1205 1645
rect 1165 1515 1175 1635
rect 1195 1515 1205 1635
rect 1165 1505 1205 1515
rect 1275 1635 1315 1645
rect 1275 1515 1285 1635
rect 1305 1515 1315 1635
rect 1275 1505 1315 1515
rect 1385 1635 1525 1645
rect 1385 1515 1395 1635
rect 1415 1515 1445 1635
rect 1465 1515 1495 1635
rect 1515 1515 1525 1635
rect 505 1455 515 1475
rect 535 1455 545 1475
rect 505 1445 545 1455
rect 450 1420 490 1430
rect 450 1400 460 1420
rect 480 1400 490 1420
rect 450 1365 490 1400
rect 450 1345 460 1365
rect 480 1345 490 1365
rect 450 1335 490 1345
rect 510 1315 540 1445
rect 560 1420 600 1430
rect 560 1400 570 1420
rect 590 1400 600 1420
rect 560 1365 600 1400
rect 560 1345 570 1365
rect 590 1345 600 1365
rect 560 1335 600 1345
rect 620 1315 650 1505
rect 670 1480 710 1485
rect 670 1475 815 1480
rect 670 1455 680 1475
rect 700 1455 815 1475
rect 670 1450 815 1455
rect 670 1445 710 1450
rect 175 1185 185 1305
rect 205 1185 215 1305
rect 175 1175 215 1185
rect 285 1305 325 1315
rect 285 1185 295 1305
rect 315 1185 325 1305
rect 285 1175 325 1185
rect 395 1305 435 1315
rect 395 1185 405 1305
rect 425 1185 435 1305
rect 395 1175 435 1185
rect 505 1305 545 1315
rect 505 1185 515 1305
rect 535 1185 545 1305
rect 505 1175 545 1185
rect 615 1305 655 1315
rect 615 1185 625 1305
rect 645 1185 655 1305
rect 615 1175 655 1185
rect 725 1305 765 1315
rect 725 1185 735 1305
rect 755 1185 765 1305
rect 725 1175 765 1185
rect 70 875 100 1175
rect 180 1095 210 1175
rect 230 1145 270 1155
rect 230 1125 240 1145
rect 260 1125 270 1145
rect 230 1115 270 1125
rect 290 1095 320 1175
rect 670 1150 710 1155
rect 565 1145 710 1150
rect 565 1125 680 1145
rect 700 1125 710 1145
rect 565 1120 710 1125
rect 120 1085 160 1095
rect 120 1065 130 1085
rect 150 1065 160 1085
rect 180 1065 265 1095
rect 120 1055 160 1065
rect 125 1030 155 1055
rect 235 1030 265 1065
rect 285 1085 325 1095
rect 285 1065 295 1085
rect 315 1065 325 1085
rect 285 1055 325 1065
rect 125 1000 210 1030
rect 235 1000 320 1030
rect 65 865 105 875
rect 65 845 75 865
rect 95 845 105 865
rect 65 835 105 845
rect 65 645 105 655
rect 65 625 75 645
rect 95 625 105 645
rect -95 525 -5 535
rect -95 405 -85 525
rect -65 405 -35 525
rect -15 405 -5 525
rect -95 270 -5 405
rect 65 525 105 625
rect 180 535 210 1000
rect 230 580 270 590
rect 230 560 240 580
rect 260 560 270 580
rect 230 550 270 560
rect 290 535 320 1000
rect 565 765 595 1120
rect 670 1115 710 1120
rect 730 1095 760 1175
rect 620 1065 760 1095
rect 785 1090 815 1450
rect 840 1150 870 1505
rect 890 1475 930 1485
rect 890 1455 900 1475
rect 920 1455 930 1475
rect 890 1445 930 1455
rect 950 1370 980 1505
rect 895 1340 980 1370
rect 1060 1370 1090 1505
rect 1110 1420 1150 1430
rect 1110 1400 1120 1420
rect 1140 1400 1150 1420
rect 1110 1390 1150 1400
rect 1060 1340 1145 1370
rect 835 1140 875 1150
rect 835 1120 845 1140
rect 865 1120 875 1140
rect 835 1110 875 1120
rect 560 755 600 765
rect 560 735 570 755
rect 590 735 600 755
rect 560 725 600 735
rect 620 655 650 1065
rect 785 1060 870 1090
rect 725 1030 765 1040
rect 725 1010 735 1030
rect 755 1010 765 1030
rect 725 1000 765 1010
rect 670 975 710 985
rect 670 955 680 975
rect 700 955 710 975
rect 670 945 710 955
rect 615 645 655 655
rect 615 625 625 645
rect 645 625 655 645
rect 615 615 655 625
rect 675 590 705 945
rect 670 580 710 590
rect 670 560 680 580
rect 700 560 710 580
rect 670 550 710 560
rect 730 535 760 1000
rect 840 985 870 1060
rect 835 975 875 985
rect 835 955 845 975
rect 865 955 875 975
rect 835 945 875 955
rect 895 930 925 1340
rect 945 1305 985 1315
rect 945 1185 955 1305
rect 975 1185 985 1305
rect 945 1175 985 1185
rect 1055 1305 1095 1315
rect 1055 1185 1065 1305
rect 1085 1185 1095 1305
rect 1055 1175 1095 1185
rect 950 1150 980 1175
rect 1000 1150 1040 1155
rect 950 1145 1040 1150
rect 950 1125 1010 1145
rect 1030 1125 1040 1145
rect 950 1120 1040 1125
rect 890 920 930 930
rect 890 900 900 920
rect 920 900 930 920
rect 890 890 930 900
rect 835 865 875 875
rect 835 845 845 865
rect 865 845 875 865
rect 835 835 875 845
rect 780 755 820 765
rect 780 735 790 755
rect 810 735 820 755
rect 780 725 820 735
rect 65 405 75 525
rect 95 405 105 525
rect 65 395 105 405
rect 175 525 215 535
rect 175 405 185 525
rect 205 405 215 525
rect 175 325 215 405
rect 285 525 325 535
rect 285 405 295 525
rect 315 405 325 525
rect 285 395 325 405
rect 395 525 435 535
rect 395 405 405 525
rect 425 405 435 525
rect 395 395 435 405
rect 505 525 545 535
rect 505 405 515 525
rect 535 405 545 525
rect 505 395 545 405
rect 615 525 655 535
rect 615 405 625 525
rect 645 405 655 525
rect 615 395 655 405
rect 725 525 765 535
rect 725 405 735 525
rect 755 405 765 525
rect 725 395 765 405
rect 120 315 270 325
rect 120 295 130 315
rect 150 295 185 315
rect 205 295 240 315
rect 260 295 270 315
rect 120 285 270 295
rect 340 315 380 325
rect 340 295 350 315
rect 370 295 380 315
rect 340 285 380 295
rect -95 260 50 270
rect 400 265 430 395
rect 450 370 490 380
rect 450 350 460 370
rect 480 350 490 370
rect 450 315 490 350
rect 450 295 460 315
rect 480 295 490 315
rect 450 285 490 295
rect 510 270 540 395
rect 560 370 600 380
rect 560 350 570 370
rect 590 350 600 370
rect 560 315 600 350
rect 560 295 570 315
rect 590 295 600 315
rect 560 285 600 295
rect -95 240 20 260
rect 40 240 50 260
rect -95 230 50 240
rect 175 235 430 265
rect -95 205 -5 230
rect -95 85 -85 205
rect -65 85 -35 205
rect -15 85 -5 205
rect -95 75 -5 85
rect 65 205 105 215
rect 65 85 75 205
rect 95 85 105 205
rect -155 30 -145 50
rect -125 30 -115 50
rect -155 20 -115 30
rect 65 50 105 85
rect 175 205 215 235
rect 395 215 430 235
rect 505 260 545 270
rect 505 240 515 260
rect 535 240 545 260
rect 175 85 185 205
rect 205 85 215 205
rect 175 75 215 85
rect 285 205 325 215
rect 285 85 295 205
rect 315 85 325 205
rect 65 30 75 50
rect 95 30 105 50
rect 65 20 105 30
rect 285 50 325 85
rect 395 205 435 215
rect 395 85 405 205
rect 425 85 435 205
rect 395 75 435 85
rect 505 205 545 240
rect 620 215 650 395
rect 670 265 710 270
rect 785 265 815 725
rect 670 260 815 265
rect 670 240 680 260
rect 700 240 815 260
rect 670 235 815 240
rect 670 230 710 235
rect 840 215 870 835
rect 895 375 925 890
rect 950 585 980 1120
rect 1000 1115 1040 1120
rect 1000 1085 1040 1095
rect 1000 1065 1010 1085
rect 1030 1065 1040 1085
rect 1000 1055 1040 1065
rect 1005 710 1035 1055
rect 1060 875 1090 1175
rect 1115 1040 1145 1340
rect 1170 1315 1200 1505
rect 1280 1315 1310 1505
rect 1165 1305 1205 1315
rect 1165 1185 1175 1305
rect 1195 1185 1205 1305
rect 1165 1175 1205 1185
rect 1275 1305 1315 1315
rect 1275 1185 1285 1305
rect 1305 1185 1315 1305
rect 1275 1175 1315 1185
rect 1385 1305 1525 1515
rect 1595 1635 1635 1645
rect 1595 1515 1605 1635
rect 1625 1515 1635 1635
rect 1595 1505 1635 1515
rect 1705 1635 1745 1645
rect 1705 1515 1715 1635
rect 1735 1515 1745 1635
rect 1705 1505 1745 1515
rect 1815 1635 1855 1645
rect 1815 1515 1825 1635
rect 1845 1515 1855 1635
rect 1815 1505 1855 1515
rect 1925 1635 1965 1645
rect 1925 1515 1935 1635
rect 1955 1515 1965 1635
rect 2145 1635 2185 1645
rect 2145 1535 2155 1635
rect 1925 1505 1965 1515
rect 2040 1515 2155 1535
rect 2175 1515 2185 1635
rect 2040 1505 2185 1515
rect 2255 1635 2295 1645
rect 2255 1515 2265 1635
rect 2285 1515 2295 1635
rect 2255 1505 2295 1515
rect 2365 1635 2405 1645
rect 2365 1515 2375 1635
rect 2395 1515 2405 1635
rect 1600 1315 1630 1505
rect 1710 1315 1740 1505
rect 1760 1420 1800 1430
rect 1760 1400 1770 1420
rect 1790 1400 1800 1420
rect 1760 1390 1800 1400
rect 1820 1370 1850 1505
rect 1765 1340 1850 1370
rect 1930 1370 1960 1505
rect 1980 1475 2020 1485
rect 1980 1455 1990 1475
rect 2010 1455 2020 1475
rect 1980 1445 2020 1455
rect 1930 1340 2015 1370
rect 1385 1185 1395 1305
rect 1415 1185 1445 1305
rect 1465 1185 1495 1305
rect 1515 1185 1525 1305
rect 1385 1175 1525 1185
rect 1595 1305 1635 1315
rect 1595 1185 1605 1305
rect 1625 1185 1635 1305
rect 1595 1175 1635 1185
rect 1705 1305 1745 1315
rect 1705 1185 1715 1305
rect 1735 1185 1745 1305
rect 1705 1175 1745 1185
rect 1220 1145 1260 1155
rect 1220 1125 1230 1145
rect 1250 1125 1260 1145
rect 1220 1115 1260 1125
rect 1110 1030 1150 1040
rect 1110 1010 1120 1030
rect 1140 1010 1150 1030
rect 1110 1000 1150 1010
rect 1225 930 1255 1115
rect 1220 920 1260 930
rect 1220 900 1230 920
rect 1250 900 1260 920
rect 1220 890 1260 900
rect 1055 865 1095 875
rect 1055 845 1065 865
rect 1085 845 1095 865
rect 1055 835 1095 845
rect 1280 820 1310 1175
rect 1330 1145 1370 1155
rect 1330 1125 1340 1145
rect 1360 1125 1370 1145
rect 1330 1115 1370 1125
rect 1540 1145 1580 1155
rect 1540 1125 1550 1145
rect 1570 1125 1580 1145
rect 1540 1115 1580 1125
rect 1335 930 1365 1115
rect 1385 1090 1435 1105
rect 1385 1070 1400 1090
rect 1420 1070 1435 1090
rect 1385 1055 1435 1070
rect 1330 920 1370 930
rect 1330 900 1340 920
rect 1360 900 1370 920
rect 1330 890 1370 900
rect 1390 920 1430 1055
rect 1545 930 1575 1115
rect 1390 900 1400 920
rect 1420 900 1430 920
rect 1390 890 1430 900
rect 1540 920 1580 930
rect 1540 900 1550 920
rect 1570 900 1580 920
rect 1540 890 1580 900
rect 1275 810 1315 820
rect 1275 790 1285 810
rect 1305 790 1315 810
rect 1275 780 1315 790
rect 1000 700 1040 710
rect 1000 680 1010 700
rect 1030 680 1040 700
rect 1000 670 1040 680
rect 1110 700 1150 710
rect 1110 680 1120 700
rect 1140 680 1150 700
rect 1110 670 1150 680
rect 1055 645 1095 655
rect 1055 625 1065 645
rect 1085 625 1095 645
rect 1055 615 1095 625
rect 1000 585 1040 590
rect 950 580 1040 585
rect 950 560 1010 580
rect 1030 560 1040 580
rect 950 555 1040 560
rect 950 535 980 555
rect 1000 550 1040 555
rect 1060 535 1090 615
rect 945 525 985 535
rect 945 405 955 525
rect 975 405 985 525
rect 945 395 985 405
rect 1055 525 1095 535
rect 1055 405 1065 525
rect 1085 405 1095 525
rect 1055 395 1095 405
rect 1115 375 1145 670
rect 1165 580 1260 590
rect 1165 560 1230 580
rect 1250 560 1260 580
rect 1165 550 1260 560
rect 1165 525 1205 550
rect 1280 535 1310 780
rect 1335 590 1365 890
rect 1480 810 1520 820
rect 1480 790 1490 810
rect 1510 790 1520 810
rect 1330 580 1370 590
rect 1330 560 1340 580
rect 1360 560 1370 580
rect 1330 550 1370 560
rect 1480 585 1520 790
rect 1545 590 1575 890
rect 1600 820 1630 1175
rect 1650 1145 1690 1155
rect 1650 1125 1660 1145
rect 1680 1125 1690 1145
rect 1650 1115 1690 1125
rect 1655 930 1685 1115
rect 1765 1040 1795 1340
rect 1815 1305 1855 1315
rect 1815 1185 1825 1305
rect 1845 1185 1855 1305
rect 1815 1175 1855 1185
rect 1925 1305 1965 1315
rect 1925 1185 1935 1305
rect 1955 1185 1965 1305
rect 1925 1175 1965 1185
rect 1760 1030 1800 1040
rect 1760 1010 1770 1030
rect 1790 1010 1800 1030
rect 1760 1000 1800 1010
rect 1650 920 1690 930
rect 1650 900 1660 920
rect 1680 900 1690 920
rect 1650 890 1690 900
rect 1820 875 1850 1175
rect 1870 1150 1910 1155
rect 1930 1150 1960 1175
rect 1870 1145 1960 1150
rect 1870 1125 1880 1145
rect 1900 1125 1960 1145
rect 1870 1120 1960 1125
rect 1870 1115 1910 1120
rect 1870 1085 1910 1095
rect 1870 1065 1880 1085
rect 1900 1065 1910 1085
rect 1870 1055 1910 1065
rect 1815 865 1855 875
rect 1815 845 1825 865
rect 1845 845 1855 865
rect 1815 835 1855 845
rect 1595 810 1635 820
rect 1595 790 1605 810
rect 1625 790 1635 810
rect 1595 780 1635 790
rect 1480 565 1490 585
rect 1510 565 1520 585
rect 1480 555 1520 565
rect 1540 580 1580 590
rect 1540 560 1550 580
rect 1570 560 1580 580
rect 1540 550 1580 560
rect 1600 535 1630 780
rect 1875 710 1905 1055
rect 1760 700 1800 710
rect 1760 680 1770 700
rect 1790 680 1800 700
rect 1760 670 1800 680
rect 1870 700 1910 710
rect 1870 680 1880 700
rect 1900 680 1910 700
rect 1870 670 1910 680
rect 1650 580 1745 590
rect 1650 560 1660 580
rect 1680 560 1745 580
rect 1650 550 1745 560
rect 1165 405 1175 525
rect 1195 405 1205 525
rect 1165 395 1205 405
rect 1275 525 1315 535
rect 1275 405 1285 525
rect 1305 405 1315 525
rect 1275 395 1315 405
rect 1385 525 1525 535
rect 1385 405 1395 525
rect 1415 405 1445 525
rect 1465 405 1495 525
rect 1515 405 1525 525
rect 895 345 980 375
rect 890 260 930 270
rect 890 240 900 260
rect 920 240 930 260
rect 890 230 930 240
rect 950 215 980 345
rect 1060 345 1145 375
rect 1060 215 1090 345
rect 1110 315 1150 325
rect 1110 295 1120 315
rect 1140 295 1150 315
rect 1110 285 1150 295
rect 1170 270 1200 395
rect 1165 260 1260 270
rect 1165 240 1230 260
rect 1250 240 1260 260
rect 1165 230 1260 240
rect 505 85 515 205
rect 535 85 545 205
rect 505 75 545 85
rect 615 205 655 215
rect 615 85 625 205
rect 645 85 655 205
rect 615 75 655 85
rect 725 205 870 215
rect 725 85 735 205
rect 755 185 870 205
rect 945 205 985 215
rect 755 85 765 185
rect 725 75 765 85
rect 945 85 955 205
rect 975 85 985 205
rect 945 75 985 85
rect 1055 205 1095 215
rect 1055 85 1065 205
rect 1085 85 1095 205
rect 1055 75 1095 85
rect 1165 205 1205 230
rect 1280 215 1310 395
rect 1165 85 1175 205
rect 1195 85 1205 205
rect 1165 75 1205 85
rect 1275 205 1315 215
rect 1275 85 1285 205
rect 1305 85 1315 205
rect 1275 75 1315 85
rect 1385 205 1525 405
rect 1595 525 1635 535
rect 1595 405 1605 525
rect 1625 405 1635 525
rect 1595 395 1635 405
rect 1705 525 1745 550
rect 1705 405 1715 525
rect 1735 405 1745 525
rect 1705 395 1745 405
rect 1600 215 1630 395
rect 1710 270 1740 395
rect 1765 375 1795 670
rect 1815 645 1855 655
rect 1815 625 1825 645
rect 1845 625 1855 645
rect 1815 615 1855 625
rect 1820 535 1850 615
rect 1870 585 1910 590
rect 1930 585 1960 1120
rect 1985 930 2015 1340
rect 2040 1150 2070 1505
rect 2200 1480 2240 1485
rect 2095 1475 2240 1480
rect 2095 1455 2210 1475
rect 2230 1455 2240 1475
rect 2095 1450 2240 1455
rect 2035 1140 2075 1150
rect 2035 1120 2045 1140
rect 2065 1120 2075 1140
rect 2035 1110 2075 1120
rect 2095 1090 2125 1450
rect 2200 1445 2240 1450
rect 2260 1315 2290 1505
rect 2365 1475 2405 1515
rect 2475 1635 2515 1645
rect 2475 1515 2485 1635
rect 2505 1515 2515 1635
rect 2475 1505 2515 1515
rect 2585 1635 2625 1670
rect 2805 1690 2845 1700
rect 2805 1670 2815 1690
rect 2835 1670 2845 1690
rect 2585 1515 2595 1635
rect 2615 1515 2625 1635
rect 2585 1505 2625 1515
rect 2695 1635 2735 1645
rect 2695 1515 2705 1635
rect 2725 1515 2735 1635
rect 2365 1455 2375 1475
rect 2395 1455 2405 1475
rect 2365 1445 2405 1455
rect 2480 1480 2515 1505
rect 2695 1480 2735 1515
rect 2805 1635 2845 1670
rect 3085 1690 3125 1700
rect 3085 1670 3095 1690
rect 3115 1670 3125 1690
rect 2805 1515 2815 1635
rect 2835 1515 2845 1635
rect 2805 1505 2845 1515
rect 2915 1635 3005 1645
rect 2915 1515 2925 1635
rect 2945 1515 2975 1635
rect 2995 1515 3005 1635
rect 2915 1485 3005 1515
rect 2480 1450 2735 1480
rect 2860 1475 3005 1485
rect 2860 1455 2870 1475
rect 2890 1455 3005 1475
rect 2310 1420 2350 1430
rect 2310 1400 2320 1420
rect 2340 1400 2350 1420
rect 2310 1365 2350 1400
rect 2310 1345 2320 1365
rect 2340 1345 2350 1365
rect 2310 1335 2350 1345
rect 2370 1315 2400 1445
rect 2420 1420 2460 1430
rect 2420 1400 2430 1420
rect 2450 1400 2460 1420
rect 2420 1365 2460 1400
rect 2420 1345 2430 1365
rect 2450 1345 2460 1365
rect 2420 1335 2460 1345
rect 2480 1315 2510 1450
rect 2860 1445 3005 1455
rect 2530 1420 2570 1430
rect 2530 1400 2540 1420
rect 2560 1400 2570 1420
rect 2530 1390 2570 1400
rect 2640 1420 2790 1430
rect 2640 1400 2650 1420
rect 2670 1400 2705 1420
rect 2725 1400 2760 1420
rect 2780 1400 2790 1420
rect 2640 1390 2790 1400
rect 2145 1305 2185 1315
rect 2145 1185 2155 1305
rect 2175 1185 2185 1305
rect 2145 1175 2185 1185
rect 2255 1305 2295 1315
rect 2255 1185 2265 1305
rect 2285 1185 2295 1305
rect 2255 1175 2295 1185
rect 2365 1305 2405 1315
rect 2365 1185 2375 1305
rect 2395 1185 2405 1305
rect 2365 1175 2405 1185
rect 2475 1305 2515 1315
rect 2475 1185 2485 1305
rect 2505 1185 2515 1305
rect 2475 1175 2515 1185
rect 2585 1305 2625 1315
rect 2585 1185 2595 1305
rect 2615 1185 2625 1305
rect 2585 1175 2625 1185
rect 2695 1305 2735 1390
rect 2695 1185 2705 1305
rect 2725 1185 2735 1305
rect 2695 1175 2735 1185
rect 2805 1305 2845 1315
rect 2805 1185 2815 1305
rect 2835 1185 2845 1305
rect 2805 1175 2845 1185
rect 2915 1305 3005 1445
rect 2915 1185 2925 1305
rect 2945 1185 2975 1305
rect 2995 1185 3005 1305
rect 2915 1175 3005 1185
rect 3025 1205 3065 1215
rect 3025 1185 3035 1205
rect 3055 1185 3065 1205
rect 2040 1060 2125 1090
rect 2150 1095 2180 1175
rect 2200 1150 2240 1155
rect 2200 1145 2345 1150
rect 2200 1125 2210 1145
rect 2230 1125 2345 1145
rect 2200 1120 2345 1125
rect 2200 1115 2240 1120
rect 2150 1065 2290 1095
rect 2040 985 2070 1060
rect 2145 1030 2185 1040
rect 2145 1010 2155 1030
rect 2175 1010 2185 1030
rect 2145 1000 2185 1010
rect 2035 975 2075 985
rect 2035 955 2045 975
rect 2065 955 2075 975
rect 2035 945 2075 955
rect 1980 920 2020 930
rect 1980 900 1990 920
rect 2010 900 2020 920
rect 1980 890 2020 900
rect 1870 580 1960 585
rect 1870 560 1880 580
rect 1900 560 1960 580
rect 1870 555 1960 560
rect 1870 550 1910 555
rect 1930 535 1960 555
rect 1815 525 1855 535
rect 1815 405 1825 525
rect 1845 405 1855 525
rect 1815 395 1855 405
rect 1925 525 1965 535
rect 1925 405 1935 525
rect 1955 405 1965 525
rect 1925 395 1965 405
rect 1985 375 2015 890
rect 2035 865 2075 875
rect 2035 845 2045 865
rect 2065 845 2075 865
rect 2035 835 2075 845
rect 1765 345 1850 375
rect 1760 315 1800 325
rect 1760 295 1770 315
rect 1790 295 1800 315
rect 1760 285 1800 295
rect 1650 260 1745 270
rect 1650 240 1660 260
rect 1680 240 1745 260
rect 1650 230 1745 240
rect 1385 85 1395 205
rect 1415 85 1445 205
rect 1465 85 1495 205
rect 1515 85 1525 205
rect 1385 75 1525 85
rect 1595 205 1635 215
rect 1595 85 1605 205
rect 1625 85 1635 205
rect 1595 75 1635 85
rect 1705 205 1745 230
rect 1820 215 1850 345
rect 1930 345 2015 375
rect 1930 215 1960 345
rect 1980 260 2020 270
rect 1980 240 1990 260
rect 2010 240 2020 260
rect 1980 230 2020 240
rect 2040 215 2070 835
rect 2090 755 2130 765
rect 2090 735 2100 755
rect 2120 735 2130 755
rect 2090 725 2130 735
rect 2095 265 2125 725
rect 2150 535 2180 1000
rect 2200 975 2240 985
rect 2200 955 2210 975
rect 2230 955 2240 975
rect 2200 945 2240 955
rect 2205 590 2235 945
rect 2260 655 2290 1065
rect 2315 765 2345 1120
rect 2590 1095 2620 1175
rect 2640 1145 2680 1155
rect 2640 1125 2650 1145
rect 2670 1125 2680 1145
rect 2640 1115 2680 1125
rect 2700 1095 2730 1175
rect 2585 1085 2625 1095
rect 2585 1065 2595 1085
rect 2615 1065 2625 1085
rect 2585 1055 2625 1065
rect 2645 1065 2730 1095
rect 2750 1085 2790 1095
rect 2750 1065 2760 1085
rect 2780 1065 2790 1085
rect 2645 1030 2675 1065
rect 2750 1055 2790 1065
rect 2755 1030 2785 1055
rect 2590 1000 2675 1030
rect 2700 1000 2785 1030
rect 2310 755 2350 765
rect 2310 735 2320 755
rect 2340 735 2350 755
rect 2310 725 2350 735
rect 2255 645 2295 655
rect 2255 625 2265 645
rect 2285 625 2295 645
rect 2255 615 2295 625
rect 2200 580 2240 590
rect 2200 560 2210 580
rect 2230 560 2240 580
rect 2200 550 2240 560
rect 2590 535 2620 1000
rect 2640 580 2680 590
rect 2640 560 2650 580
rect 2670 560 2680 580
rect 2640 550 2680 560
rect 2700 535 2730 1000
rect 2810 875 2840 1175
rect 2805 865 2845 875
rect 2805 845 2815 865
rect 2835 845 2845 865
rect 2805 835 2845 845
rect 2805 645 2845 655
rect 2805 625 2815 645
rect 2835 625 2845 645
rect 2145 525 2185 535
rect 2145 405 2155 525
rect 2175 405 2185 525
rect 2145 395 2185 405
rect 2255 525 2295 535
rect 2255 405 2265 525
rect 2285 405 2295 525
rect 2255 395 2295 405
rect 2365 525 2405 535
rect 2365 405 2375 525
rect 2395 405 2405 525
rect 2365 395 2405 405
rect 2475 525 2515 535
rect 2475 405 2485 525
rect 2505 405 2515 525
rect 2475 395 2515 405
rect 2585 525 2625 535
rect 2585 405 2595 525
rect 2615 405 2625 525
rect 2585 395 2625 405
rect 2695 525 2735 535
rect 2695 405 2705 525
rect 2725 405 2735 525
rect 2200 265 2240 270
rect 2095 260 2240 265
rect 2095 240 2210 260
rect 2230 240 2240 260
rect 2095 235 2240 240
rect 2200 230 2240 235
rect 2260 215 2290 395
rect 2310 370 2350 380
rect 2310 350 2320 370
rect 2340 350 2350 370
rect 2310 315 2350 350
rect 2310 295 2320 315
rect 2340 295 2350 315
rect 2310 285 2350 295
rect 2370 270 2400 395
rect 2420 370 2460 380
rect 2420 350 2430 370
rect 2450 350 2460 370
rect 2420 315 2460 350
rect 2420 295 2430 315
rect 2450 295 2460 315
rect 2420 285 2460 295
rect 2365 260 2405 270
rect 2365 240 2375 260
rect 2395 240 2405 260
rect 1705 85 1715 205
rect 1735 85 1745 205
rect 1705 75 1745 85
rect 1815 205 1855 215
rect 1815 85 1825 205
rect 1845 85 1855 205
rect 1815 75 1855 85
rect 1925 205 1965 215
rect 1925 85 1935 205
rect 1955 85 1965 205
rect 2040 205 2185 215
rect 2040 185 2155 205
rect 1925 75 1965 85
rect 2145 85 2155 185
rect 2175 85 2185 205
rect 2145 75 2185 85
rect 2255 205 2295 215
rect 2255 85 2265 205
rect 2285 85 2295 205
rect 2255 75 2295 85
rect 2365 205 2405 240
rect 2480 265 2510 395
rect 2695 325 2735 405
rect 2805 525 2845 625
rect 2805 405 2815 525
rect 2835 405 2845 525
rect 2805 395 2845 405
rect 2915 525 3005 535
rect 2915 405 2925 525
rect 2945 405 2975 525
rect 2995 405 3005 525
rect 2530 315 2570 325
rect 2530 295 2540 315
rect 2560 295 2570 315
rect 2530 285 2570 295
rect 2640 315 2790 325
rect 2640 295 2650 315
rect 2670 295 2705 315
rect 2725 295 2760 315
rect 2780 295 2790 315
rect 2640 285 2790 295
rect 2915 270 3005 405
rect 2480 235 2735 265
rect 2480 215 2515 235
rect 2365 85 2375 205
rect 2395 85 2405 205
rect 2365 75 2405 85
rect 2475 205 2515 215
rect 2475 85 2485 205
rect 2505 85 2515 205
rect 2475 75 2515 85
rect 2585 205 2625 215
rect 2585 85 2595 205
rect 2615 85 2625 205
rect 285 30 295 50
rect 315 30 325 50
rect 285 20 325 30
rect 2585 50 2625 85
rect 2695 205 2735 235
rect 2860 260 3005 270
rect 2860 240 2870 260
rect 2890 240 3005 260
rect 2860 230 3005 240
rect 2695 85 2705 205
rect 2725 85 2735 205
rect 2695 75 2735 85
rect 2805 205 2845 215
rect 2805 85 2815 205
rect 2835 85 2845 205
rect 2585 30 2595 50
rect 2615 30 2625 50
rect 2585 20 2625 30
rect 2805 50 2845 85
rect 2915 205 3005 230
rect 2915 85 2925 205
rect 2945 85 2975 205
rect 2995 85 3005 205
rect 2915 75 3005 85
rect 2805 30 2815 50
rect 2835 30 2845 50
rect 2805 20 2845 30
rect 3025 50 3065 1185
rect 3085 525 3125 1670
rect 3085 505 3095 525
rect 3115 505 3125 525
rect 3085 495 3125 505
rect 3025 30 3035 50
rect 3055 30 3065 50
rect 3025 20 3065 30
<< viali >>
rect -205 1670 -185 1690
rect 75 1670 95 1690
rect -85 1515 -65 1635
rect -35 1515 -15 1635
rect 295 1670 315 1690
rect 2595 1670 2615 1690
rect 515 1515 535 1635
rect 130 1400 150 1420
rect 185 1400 205 1420
rect 240 1400 260 1420
rect 350 1400 370 1420
rect -205 505 -185 525
rect -145 1185 -125 1205
rect -85 1185 -65 1305
rect -35 1185 -15 1305
rect 1175 1515 1195 1635
rect 1395 1515 1415 1635
rect 1445 1515 1465 1635
rect 1495 1515 1515 1635
rect 460 1400 480 1420
rect 570 1400 590 1420
rect 515 1185 535 1305
rect 240 1125 260 1145
rect 130 1065 150 1085
rect 295 1065 315 1085
rect 75 845 95 865
rect 75 625 95 645
rect -85 405 -65 525
rect -35 405 -15 525
rect 240 560 260 580
rect 900 1455 920 1475
rect 1120 1400 1140 1420
rect 845 1120 865 1140
rect 570 735 590 755
rect 735 1010 755 1030
rect 680 955 700 975
rect 625 625 645 645
rect 845 955 865 975
rect 900 900 920 920
rect 845 845 865 865
rect 790 735 810 755
rect 515 405 535 525
rect 130 295 150 315
rect 185 295 205 315
rect 240 295 260 315
rect 350 295 370 315
rect 460 295 480 315
rect 570 295 590 315
rect -85 85 -65 205
rect -35 85 -15 205
rect -145 30 -125 50
rect 75 30 95 50
rect 1010 1065 1030 1085
rect 1175 1185 1195 1305
rect 1715 1515 1735 1635
rect 2375 1515 2395 1635
rect 1770 1400 1790 1420
rect 1990 1455 2010 1475
rect 1395 1185 1415 1305
rect 1445 1185 1465 1305
rect 1495 1185 1515 1305
rect 1715 1185 1735 1305
rect 1120 1010 1140 1030
rect 1230 900 1250 920
rect 1065 845 1085 865
rect 1400 1070 1420 1090
rect 1340 900 1360 920
rect 1400 900 1420 920
rect 1550 900 1570 920
rect 1285 790 1305 810
rect 1010 680 1030 700
rect 1120 680 1140 700
rect 1065 625 1085 645
rect 1490 790 1510 810
rect 1770 1010 1790 1030
rect 1660 900 1680 920
rect 1880 1065 1900 1085
rect 1825 845 1845 865
rect 1605 790 1625 810
rect 1490 565 1510 585
rect 1770 680 1790 700
rect 1880 680 1900 700
rect 1175 405 1195 525
rect 1395 405 1415 525
rect 1445 405 1465 525
rect 1495 405 1515 525
rect 900 240 920 260
rect 1120 295 1140 315
rect 515 85 535 205
rect 1175 85 1195 205
rect 1715 405 1735 525
rect 1825 625 1845 645
rect 2045 1120 2065 1140
rect 2815 1670 2835 1690
rect 3095 1670 3115 1690
rect 2925 1515 2945 1635
rect 2975 1515 2995 1635
rect 2320 1400 2340 1420
rect 2430 1400 2450 1420
rect 2540 1400 2560 1420
rect 2650 1400 2670 1420
rect 2705 1400 2725 1420
rect 2760 1400 2780 1420
rect 2375 1185 2395 1305
rect 2925 1185 2945 1305
rect 2975 1185 2995 1305
rect 3035 1185 3055 1205
rect 2155 1010 2175 1030
rect 2045 955 2065 975
rect 1990 900 2010 920
rect 2045 845 2065 865
rect 1770 295 1790 315
rect 1395 85 1415 205
rect 1445 85 1465 205
rect 1495 85 1515 205
rect 1990 240 2010 260
rect 2100 735 2120 755
rect 2210 955 2230 975
rect 2650 1125 2670 1145
rect 2595 1065 2615 1085
rect 2760 1065 2780 1085
rect 2320 735 2340 755
rect 2265 625 2285 645
rect 2650 560 2670 580
rect 2815 845 2835 865
rect 2815 625 2835 645
rect 2375 405 2395 525
rect 2320 295 2340 315
rect 2430 295 2450 315
rect 1715 85 1735 205
rect 2925 405 2945 525
rect 2975 405 2995 525
rect 2540 295 2560 315
rect 2650 295 2670 315
rect 2705 295 2725 315
rect 2760 295 2780 315
rect 2375 85 2395 205
rect 295 30 315 50
rect 2595 30 2615 50
rect 2925 85 2945 205
rect 2975 85 2995 205
rect 2815 30 2835 50
rect 3095 505 3115 525
rect 3035 30 3055 50
<< metal1 >>
rect -215 1690 3125 1700
rect -215 1670 -205 1690
rect -185 1670 75 1690
rect 95 1670 295 1690
rect 315 1670 2595 1690
rect 2615 1670 2815 1690
rect 2835 1670 3095 1690
rect 3115 1670 3125 1690
rect -215 1660 3125 1670
rect -230 1635 3140 1645
rect -230 1515 -85 1635
rect -65 1515 -35 1635
rect -15 1515 515 1635
rect 535 1515 1175 1635
rect 1195 1515 1395 1635
rect 1415 1515 1445 1635
rect 1465 1515 1495 1635
rect 1515 1515 1715 1635
rect 1735 1515 2375 1635
rect 2395 1515 2925 1635
rect 2945 1515 2975 1635
rect 2995 1515 3140 1635
rect -230 1505 3140 1515
rect -230 1315 -5 1505
rect 890 1475 930 1505
rect 890 1455 900 1475
rect 920 1455 930 1475
rect 890 1445 930 1455
rect 1980 1475 2020 1505
rect 1980 1455 1990 1475
rect 2010 1455 2020 1475
rect 1980 1445 2020 1455
rect 120 1420 2790 1430
rect 120 1400 130 1420
rect 150 1400 185 1420
rect 205 1400 240 1420
rect 260 1400 350 1420
rect 370 1400 460 1420
rect 480 1400 570 1420
rect 590 1400 1120 1420
rect 1140 1400 1770 1420
rect 1790 1400 2320 1420
rect 2340 1400 2430 1420
rect 2450 1400 2540 1420
rect 2560 1400 2650 1420
rect 2670 1400 2705 1420
rect 2725 1400 2760 1420
rect 2780 1400 2790 1420
rect 120 1390 2790 1400
rect 2915 1315 3140 1505
rect -230 1305 3140 1315
rect -230 1205 -85 1305
rect -230 1185 -145 1205
rect -125 1185 -85 1205
rect -65 1185 -35 1305
rect -15 1185 515 1305
rect 535 1185 1175 1305
rect 1195 1185 1395 1305
rect 1415 1185 1445 1305
rect 1465 1185 1495 1305
rect 1515 1185 1715 1305
rect 1735 1185 2375 1305
rect 2395 1185 2925 1305
rect 2945 1185 2975 1305
rect 2995 1205 3140 1305
rect 2995 1185 3035 1205
rect 3055 1185 3140 1205
rect -230 1175 3140 1185
rect 230 1145 270 1175
rect 230 1125 240 1145
rect 260 1125 270 1145
rect 230 1115 270 1125
rect 835 1140 875 1150
rect 835 1120 845 1140
rect 865 1120 875 1140
rect 835 1095 875 1120
rect 2035 1140 2075 1150
rect 2035 1120 2045 1140
rect 2065 1120 2075 1140
rect 1385 1100 1435 1105
rect 120 1085 325 1095
rect 120 1065 130 1085
rect 150 1065 295 1085
rect 315 1065 325 1085
rect 120 1055 325 1065
rect 835 1085 1040 1095
rect 835 1065 1010 1085
rect 1030 1065 1040 1085
rect 835 1055 1040 1065
rect 1385 1060 1390 1100
rect 1430 1060 1435 1100
rect 2035 1095 2075 1120
rect 2640 1145 2680 1175
rect 2640 1125 2650 1145
rect 2670 1125 2680 1145
rect 2640 1115 2680 1125
rect 1385 1055 1435 1060
rect 1870 1085 2075 1095
rect 1870 1065 1880 1085
rect 1900 1065 2075 1085
rect 1870 1055 2075 1065
rect 2585 1085 2790 1095
rect 2585 1065 2595 1085
rect 2615 1065 2760 1085
rect 2780 1065 2790 1085
rect 2585 1055 2790 1065
rect -100 1030 3010 1040
rect -100 1010 735 1030
rect 755 1010 1120 1030
rect 1140 1010 1770 1030
rect 1790 1010 2155 1030
rect 2175 1010 3010 1030
rect -100 1000 3010 1010
rect -230 975 3140 985
rect -230 955 680 975
rect 700 955 845 975
rect 865 955 2045 975
rect 2065 955 2210 975
rect 2230 955 3140 975
rect -230 945 3140 955
rect -100 920 3010 930
rect -100 900 900 920
rect 920 900 1230 920
rect 1250 900 1340 920
rect 1360 900 1400 920
rect 1420 900 1550 920
rect 1570 900 1660 920
rect 1680 900 1990 920
rect 2010 900 3010 920
rect -100 890 3010 900
rect -100 865 3010 875
rect -100 845 75 865
rect 95 845 845 865
rect 865 845 1065 865
rect 1085 845 1825 865
rect 1845 845 2045 865
rect 2065 845 2815 865
rect 2835 845 3010 865
rect -100 835 3010 845
rect -230 810 3140 820
rect -230 790 1285 810
rect 1305 790 1490 810
rect 1510 790 1605 810
rect 1625 790 3140 810
rect -230 780 3140 790
rect -230 755 3140 765
rect -230 735 570 755
rect 590 735 790 755
rect 810 735 2100 755
rect 2120 735 2320 755
rect 2340 735 3140 755
rect -230 725 3140 735
rect -100 700 3010 710
rect -100 680 1010 700
rect 1030 680 1120 700
rect 1140 680 1770 700
rect 1790 680 1880 700
rect 1900 680 3010 700
rect -100 670 3010 680
rect -100 645 3010 655
rect -100 625 75 645
rect 95 625 625 645
rect 645 625 1065 645
rect 1085 625 1825 645
rect 1845 625 2265 645
rect 2285 625 2815 645
rect 2835 625 3010 645
rect -100 615 3010 625
rect 1475 595 1525 600
rect 230 580 270 590
rect 230 560 240 580
rect 260 560 270 580
rect -230 535 -5 550
rect 230 535 270 560
rect 1475 555 1480 595
rect 1520 555 1525 595
rect 1475 550 1525 555
rect 2640 580 2680 590
rect 2640 560 2650 580
rect 2670 560 2680 580
rect 2640 535 2680 560
rect 2915 535 3125 550
rect -230 525 3125 535
rect -230 505 -205 525
rect -185 505 -85 525
rect -230 405 -85 505
rect -65 405 -35 525
rect -15 405 515 525
rect 535 405 1175 525
rect 1195 405 1395 525
rect 1415 405 1445 525
rect 1465 405 1495 525
rect 1515 405 1715 525
rect 1735 405 2375 525
rect 2395 405 2925 525
rect 2945 405 2975 525
rect 2995 505 3095 525
rect 3115 505 3125 525
rect 2995 405 3125 505
rect -230 395 3125 405
rect -230 215 -5 395
rect 120 315 2790 325
rect 120 295 130 315
rect 150 295 185 315
rect 205 295 240 315
rect 260 295 350 315
rect 370 295 460 315
rect 480 295 570 315
rect 590 295 1120 315
rect 1140 295 1770 315
rect 1790 295 2320 315
rect 2340 295 2430 315
rect 2450 295 2540 315
rect 2560 295 2650 315
rect 2670 295 2705 315
rect 2725 295 2760 315
rect 2780 295 2790 315
rect 120 285 2790 295
rect 890 260 930 270
rect 890 240 900 260
rect 920 240 930 260
rect 890 215 930 240
rect 1980 260 2020 270
rect 1980 240 1990 260
rect 2010 240 2020 260
rect 1980 215 2020 240
rect 2915 215 3125 395
rect -230 205 3125 215
rect -230 85 -85 205
rect -65 85 -35 205
rect -15 85 515 205
rect 535 85 1175 205
rect 1195 85 1395 205
rect 1415 85 1445 205
rect 1465 85 1495 205
rect 1515 85 1715 205
rect 1735 85 2375 205
rect 2395 85 2925 205
rect 2945 85 2975 205
rect 2995 85 3125 205
rect -230 75 3125 85
rect -155 50 3065 60
rect -155 30 -145 50
rect -125 30 75 50
rect 95 30 295 50
rect 315 30 2595 50
rect 2615 30 2815 50
rect 2835 30 3035 50
rect 3055 30 3065 50
rect -155 20 3065 30
<< via1 >>
rect 1390 1090 1430 1100
rect 1390 1070 1400 1090
rect 1400 1070 1420 1090
rect 1420 1070 1430 1090
rect 1390 1060 1430 1070
rect 1480 585 1520 595
rect 1480 565 1490 585
rect 1490 565 1510 585
rect 1510 565 1520 585
rect 1480 555 1520 565
<< metal2 >>
rect 1385 1100 1435 1105
rect 1385 1060 1390 1100
rect 1430 1060 1435 1100
rect 1385 1055 1435 1060
rect 1475 595 1525 600
rect 1475 555 1480 595
rect 1520 555 1525 595
rect 1475 550 1525 555
<< via2 >>
rect 1390 1060 1430 1100
rect 1480 555 1520 595
<< metal3 >>
rect 1385 1100 1435 1105
rect 1385 1060 1390 1100
rect 1430 1060 1435 1100
rect 1385 1055 1435 1060
rect 1475 595 1525 600
rect 1475 555 1480 595
rect 1520 555 1525 595
rect 1475 5 1525 555
rect 1065 -1225 3095 5
<< via3 >>
rect 1390 1060 1430 1100
<< mimcap >>
rect 1080 -20 3080 -10
rect 1080 -55 1390 -20
rect 1425 -55 3080 -20
rect 1080 -1210 3080 -55
<< mimcapcontact >>
rect 1390 -55 1425 -20
<< metal4 >>
rect 1385 1100 1435 1105
rect 1385 1060 1390 1100
rect 1430 1060 1435 1100
rect 1385 -20 1435 1060
rect 1385 -55 1390 -20
rect 1425 -55 1435 -20
rect 1385 -60 1435 -55
<< labels >>
rlabel metal1 -230 1175 -215 1645 7 vdd
port 4 w
rlabel pdiff 830 1170 880 1320 1 net14
rlabel pdiff 830 1500 880 1650 1 net13
rlabel pdiff 2030 1500 2080 1650 1 net22
rlabel locali 1055 1505 1095 1645 1 net3
rlabel locali 1055 1175 1095 1315 1 net4
rlabel locali 945 1175 985 1315 1 net5
rlabel locali 945 1505 985 1645 1 net2
rlabel metal1 120 1390 160 1430 7 net10
rlabel locali 175 1505 215 1645 1 net12
rlabel locali 615 1505 655 1645 5 net11
rlabel metal1 -230 945 -215 985 7 v1
port 1 w
rlabel metal1 -230 725 -215 765 7 v2
port 2 w
rlabel metal1 -230 780 -215 820 7 vout
port 3 w
rlabel metal1 -230 75 -215 550 7 gnd
port 5 w
rlabel ndiff 830 70 880 220 5 net16
rlabel ndiff 830 390 880 540 5 net15
rlabel locali 1055 395 1095 535 5 net7
rlabel locali 1055 75 1095 215 5 net6
rlabel metal1 120 285 160 325 7 net9
rlabel locali 175 75 215 215 5 net1
rlabel locali 615 395 655 535 1 net8
rlabel metal1 3125 780 3140 820 3 vout
port 3 w
rlabel metal1 3125 945 3140 985 3 v1
port 1 w
rlabel metal1 3125 725 3140 765 3 v2
<< end >>
