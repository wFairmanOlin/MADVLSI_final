magic
tech sky130A
timestamp 1620813221
<< locali >>
rect 635 2090 705 2315
rect -25 1700 -5 1745
rect -85 1680 -5 1700
rect 685 1710 705 2090
rect 5730 2090 5800 2315
rect 6470 2090 6535 2315
rect 685 1690 3410 1710
rect -25 1020 -5 1680
rect 3390 1630 3410 1690
rect 5730 1630 5750 2090
rect 6515 1710 6535 2090
rect 6515 1690 9240 1710
rect 9220 1650 9240 1690
rect 9220 1630 11450 1650
rect 3390 1610 5750 1630
rect -45 725 -5 1020
rect -45 705 -35 725
rect -15 705 -5 725
rect -45 695 -5 705
rect 5730 730 5750 1610
rect 5730 720 5770 730
rect 5730 700 5740 720
rect 5760 700 5770 720
rect 5730 690 5770 700
rect 5655 425 5695 435
rect -145 365 -45 415
rect 5655 405 5665 425
rect 5685 405 5695 425
rect 5655 395 5695 405
rect 11430 430 11450 1630
rect 11430 420 11470 430
rect 11430 400 11440 420
rect 11460 400 11470 420
rect 11430 390 11470 400
rect -80 -840 -45 365
rect 5655 335 5695 345
rect 5655 315 5665 335
rect 5685 315 5695 335
rect 5655 305 5695 315
rect 5675 245 5695 305
rect 5365 225 5695 245
rect -80 -850 -40 -840
rect -80 -870 -70 -850
rect -50 -870 -40 -850
rect -80 -880 -40 -870
rect 5365 -1745 5385 225
rect 5730 -845 5770 -835
rect 5730 -865 5740 -845
rect 5760 -865 5770 -845
rect 5730 -875 5770 -865
rect 5655 -1370 5695 -1360
rect 5655 -1390 5665 -1370
rect 5685 -1390 5695 -1370
rect 5655 -1400 5695 -1390
rect 5750 -1755 5770 -875
rect 5710 -1780 5770 -1755
<< viali >>
rect -35 705 -15 725
rect 5740 700 5760 720
rect 5665 405 5685 425
rect 11440 400 11460 420
rect 5665 315 5685 335
rect -70 -870 -50 -850
rect 5740 -865 5760 -845
rect 5665 -1390 5685 -1370
<< metal1 >>
rect -110 1050 40 1085
rect 0 955 40 1050
rect 5470 910 5795 950
rect -45 725 15 735
rect -45 705 -35 725
rect -15 705 15 725
rect -45 695 15 705
rect 5470 345 5510 910
rect 5730 720 5795 730
rect 5730 700 5740 720
rect 5760 700 5795 720
rect 5730 690 5795 700
rect 5655 425 5695 435
rect 5655 405 5665 425
rect 5685 405 5695 425
rect 5655 395 5695 405
rect 11430 420 11470 430
rect 11430 400 11440 420
rect 11460 400 11470 420
rect 11430 390 11470 400
rect 5655 335 5695 345
rect 5655 315 5665 335
rect 5685 315 5695 335
rect 5655 305 5695 315
rect -80 -850 0 -840
rect -80 -870 -70 -850
rect -50 -870 0 -850
rect -80 -880 0 -870
rect 5730 -845 5805 -835
rect 5730 -865 5740 -845
rect 5760 -865 5805 -845
rect 5730 -875 5805 -865
rect -5 -1100 15 -1005
rect 5790 -1055 5845 -1040
rect 5655 -1370 5695 -1360
rect 5655 -1390 5665 -1370
rect 5685 -1390 5695 -1370
rect 5655 -1400 5695 -1390
rect 11430 -1395 11445 -1355
<< metal3 >>
rect 3510 1610 5475 1630
use 10k_res  10k_res_3
timestamp 1620799792
transform 0 1 5165 -1 0 -1745
box 0 0 35 605
use opamp  opamp_2 ~/Desktop/MADVLSI_final/layout
timestamp 1620660520
transform 1 0 230 0 1 -1825
box -230 30 5425 1700
use 10k_res  10k_res_2
timestamp 1620799792
transform 1 0 5695 0 1 -1400
box 0 0 35 605
use opamp  opamp_3
timestamp 1620660520
transform 1 0 6020 0 1 -1820
box -230 30 5425 1700
use opamp  opamp_0
timestamp 1620660520
transform 1 0 230 0 1 -30
box -230 30 5425 1700
use 10k_res  10k_res_1
timestamp 1620799792
transform 1 0 -80 0 1 415
box 0 0 35 605
use 10k_res  10k_res_0
timestamp 1620799792
transform 1 0 5695 0 1 395
box 0 0 35 605
use opamp  opamp_1
timestamp 1620660520
transform 1 0 6020 0 1 -35
box -230 30 5425 1700
use 50k_res  50k_res_0
timestamp 1620810761
transform -1 0 630 0 1 1705
box -5 -5 670 610
use 50k_res  50k_res_1
timestamp 1620810761
transform 1 0 5805 0 1 1705
box -5 -5 670 610
<< labels >>
rlabel locali 11470 410 11470 410 3 Vint
port 1 e
rlabel metal1 11445 -1375 11445 -1375 3 Vprop
port 2 e
rlabel locali -145 385 -145 385 7 Verror
port 3 w
rlabel metal1 -110 1065 -110 1065 7 Vref
port 4 w
rlabel locali -85 1690 -85 1690 7 Cap1
port 5 w
rlabel locali 700 2315 700 2315 1 Cap2
port 6 n
<< end >>
