magic
tech sky130A
timestamp 1620757311
<< xpolycontact >>
rect 0 385 35 605
rect 0 0 35 220
<< xpolyres >>
rect 0 220 35 385
<< end >>
