magic
tech sky130A
timestamp 1620530725
<< metal3 >>
rect -15 -15 1015 1015
rect 90 -45 135 -15
<< mimcap >>
rect 0 45 1000 1000
rect 0 10 10 45
rect 45 10 1000 45
rect 0 0 1000 10
<< mimcapcontact >>
rect 10 10 45 45
<< metal4 >>
rect 5 45 50 50
rect 5 10 10 45
rect 45 10 50 45
rect 5 -45 50 10
<< labels >>
rlabel metal4 25 -45 25 -45 5 top
rlabel metal3 110 -45 110 -45 5 bot
<< end >>
